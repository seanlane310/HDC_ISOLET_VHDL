library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
 
entity testing is
end testing;
 
architecture behave of testing is
 

	type slv_arrayclass is array (0 to 5) of std_logic_vector(9999 downto 0); -- length of this array must be number of classes (letters) we are tested, vector length is dimensions used
	type testarray is array (0 to 5) of std_logic_vector(9999 downto 0); --length of this array must be number of test inputs we are running
	type testactual is array (0 to 5) of integer; --length of this array must be number of test inputs we are running
	type samearray is array (0 to 5) of integer; --length of this array must be number of classes we are using
  	signal result : integer;
  	--signal total : integer;
  	--signal correct : integer;

  function classification(
    testinput : in std_logic_vector(9999 downto 0);
    classes : in slv_arrayclass)
    return integer is
    variable closest: integer:= 0;
    variable mostsame: integer:= 0;
    variable numclasses: integer:= 6; --number of classes (letters) we are checking
    variable numdimensions: integer:= 10000; --number of dimensions for HVs
    variable same: std_logic;
    variable amountsame : samearray := (0, 0, 0, 0, 0, 0); 
  begin

  	L1: for i in 0 to numclasses-1 loop
		L2: for j in 0 to numdimensions-1 loop
  			same := testinput(j) xnor classes(i)(j);
			if (same = '1') then
				amountsame(i) := amountsame(i) + 1;
			end if;
		end loop L2;
		if (amountsame(i) > mostsame) then
			mostsame := amountsame(i);
			closest := i;	
		end if;
  	end loop L1;
    return closest;
  end; 
   
begin
 
  process is
-- store classes in test class array 
-- store test inputs in test as an array of test inputs
-- store the actual value of the test (whether a,b,c,etc.) in testactual array
-- store number of tests you are conducting in numtests
-- loop will run tests with each of test inputs to find what class it most closely matches
-- it will return that index as result
-- if index matches the actual expected result index, correct counter is incremented
-- the total number of tests conducted is incremented regardless of correct or incorrect prediction
 	variable testclasses : slv_arrayclass := ("0001010001010110001000000100100011010111100000011100011000100100000011100000001010000101010101000000101100010000001100100000001101000111111001111000011010010010000100001100100000011001000001000011010000000001001000001000100101010100100000100000001000100010010100000001100000000100001000100000011101100011001101001100010000000000000111100000000100001000000010110000001100000000110000001010000000001010010000111011000010110000000000000100001001010100011000000100110001001000111000100000000010100101100000101000000000001000000000000000000000010000110000000100101100010001001100000001000100000010110100000000000000110000001110111000000000010001000100000000000010000001111000110000010000000001001000000000000010000000000000011011001100000010111001000010000000101000110000000100110000100010001000000001000101000001001000111100000101010000000010010101000100000010000011000110000000000000010001100000001001100010001000001100000000110000000100100001011000101000001100100001110010101100000110001011011000110100100001001100000000110101001001111000001011001110000001000010101000000000100101010000000000011001010000110010001001010000010100010000001001111000001010000000000000100000010110000011000010100001101010100100010010100101101000001010010000000010010000000010011000000000000000000110000110101100101011001000010100100100000011010001010000101001000100000010010001000010000000001001010000010001000100100000000100000001000000010000110100100010000000001010100000000010010001110001000000010000000000100000010000011100010001000000010000100000000000001000110010001000011100111000110010000000001000010000101010011010000000100111000011000000101000000011011000011000110000010000100000000000110000100000000000000000000000100110100100001100011000101000000000000010000000000000000000101001000001011010000001001010001000000001010110100110010010010100000001000010100101000001100100000100001001100011011000011000100000010010000000000010010100000110100101000000000000000110011010000000000001011000000001000000000001010001000000000000000000100001100000110001100001001010000001100100000000100010100000100100100010110001010100100000000001000000000000001010000001000100010001011010000000000100100000011000001000011000010010100000100001100001010010010000010000010000010000100000111001000010000000100000110010000100010000000001000010100001010010001000110001110100000111000101010010000001010000000001010010010001101011111101100001100001000000100000000000011001100010001000000000010000000000000100000100100000110000100000000000011000000010000000101101000000100100100110000000101010100000000000100000010000000001000000101110000011000000101101010001100100010000000000110001001001000101000100000000101000000100011000111000010000001001010000010101010100010000000001001000111100000111000100001000001010001000100111100000000000010000000000100000001001000100000000000000010000000000100100000100000000100100011000010001000001001000000000001000100011101000010100010000001010101101000110100000010000000000000100000101000010000000101000000000000000101000111110000001000000000000001000000000000101011100110100011000010000000000000010000000001101100000010000101000000010000100000101101100010000001010000000000110000100101100100010000001011010001000000001001100100000010100010100100000000100101000000001001001011100010001000100000000000100000000101111000000000000000100101000000010000000100001000001101010000100010001001001110000001000011000000100100000000000010000010111000100100010000000000100000010000011000100100011100101000000001011010000001000101000100010010000100001010000010010010000100000011100001001011100100000011010000000100000000111000001010100101100101100000001100000000011000001000000100010010001010010010100010111000000010000010000001100001101000001100010000110000000100101000000000001000101100000001110100100010000000100000000000010000000001000000000010000011010000000001101010000000110000001001010000100101000000000011000000010001001000000001000000010000010111100100000000011001001000000000000000010000001001101000010011000000100010000001100000110000001100110100000010000001000010000000001000010110000101101001000001000000101000000011000000000000010000110010000010000001000000000001000010000011000000000000000010011000000001100010101000101000000111001000000000000000011010000001010000110000000001000101001110010010000100001000000000000010000000001000000000000000010000100000000100000001001000100010010010001000100000000000011010010000110010000100100010100001001110000000000001000110010001110000000000000000001100000000000000001011000000000110000100001110101000000000001000100100100000110000010000100000100010101000001000110000001010000000000010000000000001000010100000011000000000110110010100101000010001000111000001100010011101110001100011000100001000000100100000000001000001000000000010011000011011100010001001000000100010010010000010000110010100001000010000000010111010011000101000000110100001000000000010000010011000000101001000000100100000000001000000000000000000000101000000101011000000000101000000001000111100100010000100110000100010000000000000001001000010010000000000000000000001000000010100010000000001000011000000111110101101000100101100011000000010000000001110110100100010010000101000000001000000100000110000100000000000100001100000000100010000100000100010000010110101100000000011011000100001000010011000000000000000000100001000100000000000011010000010000001000001000001011000001000100000010000011100000101100001000010100010111100010011100100010000001000010000000100000100000000000100000010010010100000100100110000000000100000101000000001100010000000000000000000011000001010000000100000010101101000011110001011000000101100011100100000000010000000010000000000000000100000000000000010101000010000000010000000010110001000011100000000001100010100101000110100001001000000101011000000000000000000001001000100000110000010101011000000000101010000000000110000001011100010000010001010000111010000100000110000000010110000000000011100100100011100000010000000000100000001101101000000000000000110100100100000001101000010101010100001000000000000001000010111111001000010100001000000000100100001110100000100000000101000000011110100000001010001100001011001000000000001000000000001000000000010000000001000001000000000110010010000000011000001001000001000000110000001000010000000000001000110100010001000000110000011000011000001100010010001000001001110100000001100010000010100000000100000001001000001000000011011000000100010001000000001000001000000000001100000000000000110000000000100100010000001000000000100001000011000000011000000100000100001000100010010000000100100010000100100110000000010010001110000001000110000110010110110000011000000000100000000010100011000000000000100001110000000010000110000000010000110100000001000100010101000000000000000000000000011100011000000000100100001100000110001100101000001101110000011010000001000001010001010000100000000000000100000000000100100011101010000000011000010000001001001110000010000000000000010000100000010000100110000000001010010000000110010000001010000100001000100100000010100000000000000000101011010001001000000001000000011000001000101110000000000001001001000000100010111010000010001000110101000001110011111000100000001000001011000110000110100010000000000000000010110011000001100000000000000100010000111101100010000000100001010000010001000001000000000110100110101101110010100000000011001000001001000001000100000100010011101001001000010010000100100011100000000000000010001000110000000100100100100101010110000111010000101000010000000100000000000101000000111010000100100000001000000000011100001010000011111111010001001000001001000101000010000100000000011100100100000000010000000000000000111000001000011011000000000000000101000010101000000000000011110010001101000001101001010001010000010001010000100110101011101100000111011101001010000000100100010000001100101010000010000000010000001100100011000000010000110001000000111000000101111000000001000000000010000000100001000001000000000000000000000000000000100000100000101000100000000000001010110000111000000000010000000000000000010000001000101011000100000000000100001010010100000001001100010000000010000111000110100000001001011010000010100101011000000001000001000000010010000010100000000100010000000010001101001100010010111010100010100010000100001000000010000010000000000001000001000011001010110010000010000000010111000100100000110100110000001000000010000011000000101010000110000000100100011110101110100000000000100010000000101000100000000010000000011000010000001001000000001000011000100000000001000000000100100011000010010000100111000100100000000110010010000100000000001010001000101001000000000000100000001100010001000000000110000000110001001000000100110000011101000000001000000000001110101000100000010110000001000101000100000000001100110100000101001101011110010000001100000000001100001000010001001000011001000001011100110010100000001000100001000000001011000000000111011000001000000000010000000011001000000011010001101000100010000110100011010000100001001010001000101110100100100000000100000100001011000000000000001001100000010001000001111000000000000000000100000000000000010001000000000010100000000000000000000010010000011000000100010100000000010000010001001010000000011000000000001000010000000000100011000001010011100001000000001100001101110001000000000010000100000010001011100100000000010010000100000110010001000001100000000000110000000011100000000001101010000001100101100000000110010000000001000100000000010101000000000000000100000000100010000000000001000001000100000100010001010011000100100001001001000000100011000011010000101000001110001011000000000010011000001011100010000000000000001100010001000101000010100001001000100001010111001010111000101100010000010000101000101000010001101001000010110000101000000100000001111100100001001100010101100000000000000001000110100100001010000001001100011100001000010000001000001000000000010000100000000110110000110010011111000010001110110101000010100101000001001100001001010000000010101001000100000000000010000000000010101010010000100100001001010000000000000001000000000001011000000010000100000100000011010110",
	"1011010001000000100000000100100001110100100000010100010001000100100010100000000010001100000101000100010110011000100100100010000111100001110000111000011010010001000110000000000010001101010000000010000000000001001000001000000101000110001000100001001000100000010000000001101000000101110000100000011100010101001100001100010000000000000101100001001000001000000000111000000100100000110001001000000000001110001000001000000000110110110010010001101101010100000000001000100001001000101001000100000000000101100000101000000000000000000000000000000000010000001100000000000100010001001001000001000110000010110100001000010000000001000111010000000000000011010101010001000010000101111000000010000000001000101010000100001110100000010000001011000100000000101101001010010000101000111000000100000001001000001010000010000111010001101000010100000101011100010011000101000010001011000001100110000101000010010000100000001010110011010000001100000000110001100100100000011000111010000100100101100010000001100111101000011000011101000000001101100000110100001001110000001101000110100001000010101001011001000101010000100000000000011010111010001001000000010100010000001101110000000100000001100000100000010111000101000000100000100010000111110110000000000011101000010000001010010000100011000000001000000000000100000110011001101010001000110100100110000011000011010000001101000100000010000001010010000000000001000000000001000001100000001100100000001000010000110000100000000000000010100000000100011001001001000001000000000001100100110000011100010011001001001000000100000000001000111010001000101100011000111010000010101010010000011000011000000010000111100011010000100111100010001000011000110100010001000000010000100100101010100000100000100000010100000001000110101001100101100100000000100100000000000001111011000000011010000001010010000000001001010100000100011000001100100100000010010001001001100100000000001001100010010000010101010000001010100100100010000110000001101000001000001000000110011010000000000010011000000001000000000000010001000000000000001000000100100100010001000111001000000001100110000100100001100000000100000010101010010100000100000100000000000000000100000010000000110000010000000001000000000000000000000000001010010011000000101001100001010010010000000001000000010100100000100001000000000000100000000010000111010010001010010110000011110010000000110000110000000110001000010000000100000100000000010010010001100110011001100011010000000000000000000000011001001010001100000001110000001000000000000011001000100000100001000100011001000110000000101000001000100111000000000000000000100000000000100100001000100000000000101110010100010001000000010001101100000000000001000001001001000111000000010000101010000100010001111000010000000001010000010001000100010000100000101000001000000010001110000000100011001000010011100000000001000000010001100110011001000000000000000100100000000000000001000100001000000110011001000001000001001000000000001000000001101000100000000010101000001101001100000100010000000010100000110101001000001110101001000000110001001100100100000001000010000100000000000100000100010101010000011000010000001001000010000000001101000010000100001000000010000100100101100100010000001001000000000000101100000100101000000000011010000001000011101000000000001000110100100000000100011000000001000001011100000100000101000000010000000100001110000001000000000000100000000010010001110101011000100010000100010001001000100001010000011000000000100100010000010000010000010000110000000000100100000010001001000000100001001000000001010001010000001000011000001000010100100000010000000000010000100000000100001001011001100000010001000000100000000010000001010100000000100000000011000010001001011000000101000011010011010000000000010101000100010000010010101010001000110001100001010011000000000101000010000001010101100001101110000100000000000100000000100010000000001100000000010000000000000010001101010000001110000001101000001100101000000001001100001100000011000010010100000000010010100100100000000011001000000000001010000010000000011100000010011000000000010010001000100110010001000100100000110000011000000001000001100000000000100000100010101000000101000000011001000000001110010100000010010000001000100001001000010000011100000000000000111000100000000101000001000101000000001000000000010000000010110000001010000110000000101011001000110000010000000000101000011001011111000011000000010000000110000100000000100000000011000001010000010000100000001000000001010000000110010001000110000000001001100001000000011011110010001110010001000001000101110100011000000001001100000000110000000000110001000010000010000000110000000110000010000000000100010001000001000010011001010000000110110000000100001000110110000000001001100110110010100001001100000000110000000100010010100010001000011001100000000000000100000000000000001000000000010001001001101110000001000100101100010000000000000100110111100001000010000010110010010011001000001000110100101010000001000001011101000000101001100000100100100000001000000000000000000010100000000101001000000000101110000101000101101100010001000100101100100001100000000011000000010000000000001010000011000010010000100010011100001001000001100110111000001000110001100011000000000000000001010100000000010010100100000000001000000100100000011000000001000100001101010000000010110101001101010000001110000100000000001001000100001000010010001010000001001000110001101100000000000001010000000000000000011000000000000000000100001000001001100000000011001000010100010101101010000000100010000001000000110001010010000000000010100010010011110000100101100010000000000001000000000000001000010000100000010110000001100001010011000100000010111001001011100001001000000001100011100110000000101000000010010011000101000000000010000000010101000000000000010000001100110000000000010000000000100010000101100010000001001100011100111000000010000000000000111010100010111000010011010000000000001010011000000110000101000011010000010000000000011000010010000110000000010010010000000010100101110010100010100000000000000000011101001000000001100110100001000100001001010000000100010010001000000010000101001110001011001010000000001000000100100001011010100000000000101101100000001111000000000010001101100101111100000000000000000000001001000000000001010000000001001000000110000010000000011001001001000100000001010000001000101000001000001000110000010000100000010000011000001010000100010000100010001000110010000001110010000000100000000101000001010000000000000011001000001100000001000000000000000000000100000000000001000000100000000000100100010000010100000000000011011011000000010001001100101100000010100110010000000110000010010010000010010001100010000100000001100100000100010110010000011000100001000011000000000101000000011000000101110000000010000110000000000000111100010001010100011101000001000000100000010000100100111010000000101000011100000110101100010000001101100000010010001000000000000011010001100000000010000000000000000100000011101101000000110000010110001001000100000010100001001000010000100000100001100110000000001010010000000100010010001110000100101000100010000010000000100010001010010000010000001000000100000000011110000001001010010000000101000010000000000000010001000010001101110100000101110010111010000010100000001011000010010010101000001001100000100000000010000000100000001001000100100000111100100010000010100001010000010000000001000000000110100100000100110000100001001011000110010001000001000101000000010111100000000000011010100000100010000000001000000010001010000010000100100001000100010100000111000000011000000000000110000000000100000100001010000100100000000100000000001110000010000010001001010001001000100001000101010010010001100000000000000100100000010000000000000000110000000000011000001000000100000011001000101000000000101011010000001010010000111110100000010000000010010001010010001010001000000100011001000000101000101100010000001000100010000010001100011000101100000010000110010000010110000000010001000001111000100011000000000010000000000001001001000000100000001100000000010010100000100000001000100000001000001010100000100100000000000100000001010110000001111000100001001100000001010010001010001110000101001000000100000000000100100001100000110001010000000110100100000000000001000001000000010010010000000001000101010000100010000100000000000010100000000010010000100101000000011010000110011000000000000001000001001010111010000010101000010111000000100010110100100000000000010000110011000000100010000110100000101101011010111000100000000000100010000011000000011100000000101010111000000000001000000001000101001100110000000000100001000100101001100000010010110110000100100010000100010000000100010100100010001000100101010100000000100000001100001001000100100100000000010001010000000100110100001100000000001000000010100110110000000000010100000010100010001100000000001100100101000100010010011110010000001000000000101010001000000010111000001000000010001000110010100011011000100100010000001001000000000100000000100110000010011100000010001000000001011101011001100010001100100111001000110001100010001000101010000100100001100001001000001001100000000000001101110000000001000110101000000101000000100100000001010000010011011000000010101000001101000010110000010010011001010000000100100000010010010001000011000101011000000000000001010000110001100010011010000001100011000001100010001110100000000000000000000000000010011111000000100000010010010100000011010000100001100010000001100000100110100000000001000000000001100000100000101110010001010001010000000000000101000000000000000100000000000010001010100111000011000000000100000001010111000000000100001000000000001001000001000000100001001110001011000000000011011001001000100010000000000001000000010001000001000001100001000100010000010000001000110100000101000000010000100010100000011000101001001000100000101000100100000000011100110001101000000001000000000000000000100100001100001010000100000100011000001000000000101010001000000000000001010000001001100000110011110101000010000100100101100010010100000010000110000000000010000010001000100000100000000000000001000000100100110000000100000000000000000001010101000101000001100100000101000100000100101100010000",
	"0101010000010010001000010100100000011110000100011100001000010101100101100000001000001101010000000000101100001001001000000001011001010011011000011010011000010010100000010000100000011001000001001011000010000000001000001000000111000100101000000011000000100010010100000001101000000100101000100010110101000101001101000000010000001000001100100011001100000000000000010000011110110000010001000010001000001100011100110010000110110111010000001101101101001010001100100100100000000000111001000000000100100000101001100000000000000000010000001111000000100011000000000100000000010000001101000001000100001000110100001100010000100001001100101000000000010011000101010001000000010100011000010000000000000001101001000100001010001100000000010011000100000010011101000000100000001000110011000100110101101010000010000011000000001100100000111101000011001000011110000101001010101010000001000100000100000000110001000010000000010011011000001001000000110101100010100000000010010010000100100001010110101101100001000001011000000001000000001001000000100001000001100000001101000000000000100000101001010000011001010000001000010000000000100000001001010100010100000000011001100001001110000000000010000000000110010010000011000101100110100001000010000000110111101000110100000000010000000011011000101000000000010111111000100100001010001000000101000010000011011001010000001100000100000000000000011010000001001000010000010001000000000000000100100100100000010100010010100000001010001010110001000100010000010001000000010100000000100100110000011100110011101000000000000000100000000000111000100000101100011000011010000000001000110000111000011000100100000001000011010001001101000011011100001000100000000000100000000010000000101010000000000100100000110010000001000010001000100001000100000011000000000000010001001000000000011010000001000010000000000001010111000111010010010001000001000000110100001000100001001100011001000110001000010101001000000010100000110010011011000100000001001000001000000000001000000000000001001000000000000000101001010001000000000010000000100001101000100001000000010000000001010110001000100010100000100000000010011001000000100000010101000000000000001000000010000100100000001011100001100100101000011100101100011010010011100000100101000001100000011000000000000000010100000000011000010011000000100000100010100011000010000000010000100011010010001000110000110000000110000101000010000101110100001001000010010000001111110000000001110000000000011000000001100001000110001000000000010000001000000100000010110000011000101000001100000001000010000000101000000001100100100100100000000010100000000000101100001011100001000100001100000100000000000110010001101100000000001001100000001001000110000100010000001111000000001000111000000000001000100000010001010000000000100001100000001000000111001000110000001011000001101111000000101001010000010000100000000000000001100010000001111000000000000111000000001000101000010001000000000100000000000000000000100101111000000100001000001010001101000010100100010000100000100001010101001000000100111110000000010000101000101100000100000000000100000001001101000100000100101000010100010000000000000000000000000101100000001000001000000110000000100001000101100000000001000000100010100100001000101000000001001000001000000010001101100000010101111100101000000000001000000000000000000100010000000001000100000001000101000001000000000100000100001010010110010101110001100000011000000000011000001000100000001000001010000100100110010000010000010110000000010100010010000100000000000000000100000010100100000001001011010001001000100010101010010100000000000000001010010100100000010000000000011011000000000011000000100000000100000001000000001000100100000011110000001011011001000000000010010011010010010100010010000000000000000001101010001100110000110011000000001000101001001000000001110111000000001000000101000000001000100000000110000000001000000000010000001010100010001100010100000010010001101100000000001000000001011000001010000001000010011100000010010010100100101000010011101000100000000010000010000001011100000010000100000100010110000000000110000001100100100000000000001000000001000000000010101000100000100000100000000101100001001001000000000110010010010010000110000000000001001000010000010000000000000000110001000000100101000111000100000000011000100000000001000001110000000000000000000011000001100001010000010001100000011100010000011001000011000000010000000100001100100000000110000000000100001000010000100100000000000011000011000111000001100110000001000001100010000000001010110000101100010001000000000001100100010000010001010000000000000000000101000101000000010011000101100100010010000000000000001000000101000101000101001101010000000000010000000000011000100110000011000011000110010010000100000011000000000000000101010000001100000001111011111010000010100000011000101000010001000001000111001010001110000001001100001000010000100000010000000000100001000000010010010100010001101000011000010100100010000000010000101110100010001001110100000100100000000000100000010000000010100000000101010000010000100010000100100011000000011000010100111100010010100000011000001000000010000011000100000000000010010000000010001000001000011000000101010000101001110101100000000100000000001001000100100100010000011101010000001100000000000110010100010001000100000100010010001011010100000101011001101010111100100100011010000110001000010010000000010000011100100001110000010000000001010000100000000000001000001011000000100001000100000011100010100001000000010100000000101010010000000010000100001010110001100010000000100001000000010011010000100000100110000000000100000001001010001100000000100000001010000001100001010100101000001001101101001111110001011000000100100000100000000000100010000000000010000000000110000000000010000000000110000010110010001010010100000010100000101001100110001101011110110000000000000000001000000010010000001001010000101010111000010011010000011001101000001010001010001101001011010000110110010000110010110000110110000000010100000000001011100001010000000000111000000000000000110001100000000110100011110101100110001100101100000100010110000000000000000001001000100000001010010100000001000100000000001100100000110100101000000001010110010000001100000001000100010000000000001100000000001000010000010000000001000001101001010010011000000001010001001001000100010001100000001000000100000010001100110000000000110010110000011000011010001100010010111000011000110110000001000010010011000000000101000000011000011000000001011000001000110010000000000001001001100100000100000001000000000010000000000000000000011100000000100010000000000000000001000000000110000010100110010001000000000010000110010000010010100000000110100001100010000010010110110000010000100001100110000010000001100000001000100101110000000010010110000000000000011110000011110100010100001000010000101000001000101100011000000000100000011100000010100100001011001101010000011010001101000001010001100000000000000000001000000100000100000001101001000000001000010000001001000110110000101100001000000000101000010001000010000000000011010010000110100110001100001000100000100111000001100001000000001000001101000001001010000001100000010110000100101000000000010101001110000000000000011011000010000100000001010001000111001000000000001000000001000000010110101010000011101000001010110001000001000000001000000000010000100110100000001000100000010000010010010001000001000111000100000100100010100000100001001100111001000001000000000101010010000000000000011100000100100010000000000000100010010000110000000100100000100011110000000011010000111000000000100111000000000101000000000010000100100010001100000000000100001110000000000111010011000010101000010100010010000100100100000100101000100000010010000101001100110000001000011010001000100100100010001000101100001000001011000000000010010000011110110000010000000000010000011110001101001000000110010100000010101000001000100100000100010010000110001000000000100000100000000010010000101101010000010001100101110000100011000010000010000000000000000001010010000000001000000000100001100001100000011000000100001000001000000000110100000000000000000001010010010000101110101001000000000000000110001101001100100001001111000000100010000010100000100101001011000110000000000101101000000000000100000000000000000010000000000100010000101000101001001001011010011010100010000110000001001100111010000010011000000001000001000111000000101010100100100001000110000100000010110100010100001000000000010001001000100010000010100000100000010100100110000100011000000100100011000000011000000010000000010000100000001001000001001100010000000000000000001011001100100011000000010000000101000100000010000110001000000000010101111010100000001101000000000000100101001100010001000110100100000000110001110000000001110000010100000000100001000000011110000000100000000010010010100101010100000000011000100000000001010111000000010100000100000000100010000011001001001100001100001010000000110000100000010011000001000000001010000000000011111000101000000010010000000011001000010011011001000101000000000000100011000000000001100000001000010010000000101101100000000100000010000010000000000100010000001001000101011000010000001010100000001101010000000010010010000010000000101000000000010000010001011000000000010000100000010000010001001101001001010000100000000010010000000000110010001010010010101001000001000110101100100000000000001010000001000010011101100000000010010000010000000000010001100011110110001001100100000111000000000001101011000001010101000000000000000001000100001000001000110101000000000000000100000000000000001010110011100010000010010000000001000000000100100101001011000000101001000011110000001000001100000001000000001001001000001010010000000000000100000110000000000101100010110001001000110000010101101010010100000101000010010000001000001010000001100000000000010010101000000100010000101100101000000000000101111000000001000000100110000000001010000101001100011100000000010100100100001000000000000000100000001111110000010010100111000010001110000000001000100001101011000010000000110000100010000001010100011010000011001000000110101100100001100000000001010010100000010000000100110001000001100100000000000111101010100000",
	"1001010001010100001000000100000000011111100001011100011000010100000011100000001010001001000001100100101110001000001100100001001011100011011001011000001010000010100000000100100001011001000001000011000000000000001000001000100101010100101001000001001100001000000000000001001000000001001000100001111000001111000001000110010000001000001110100011000100001000000000110000011110100000110000001010001000001100010100100001000100010110010000000000000000010101010000001000110001001000101001000100000110000100001001001000000000001000011010100100000000011000101000000000101000010000001000000001000100001010110100000100010000000001001111011000100000010000001000000000000010011001100000110010010000001001101101100100001110001000010000001011001000000010010001001011000000101000111010000000010101100010011010000001000011001000000000111101000000001100000110000101000000000011000011100110000000000010010000000000001010100001001000000001000100100001000000100001010010110000001100100101010010101000000101100010011000111101100001001101101000100001001000100001011101011110000011000010000000011000001100010000101100011001010000010000001000000010010100010000001101001000010101000000001000100000010111010101000010100001101110100101110000000101011011001010110100000000010000100010010000101000010000010101000110101100101011001000010101000010000011011001000000101000000100010010000001011010000001000000010000000001000000100000000000010000100000010000110000100010000000000000110001000000011100011001000000010000000001100100100000010100110010001000011010000001000000000010100000001000101100110000111010000000001000110010000010001000100010100101010111010001001010100011011100001000100100010000000000000000100000101010100000000000100000100010100101001010011001100100000100000001000100000000000011001001000000011000001001001010000000000000000100100011011010010100101000000000100101001001110001001100001001100110011000011000100000111010100100100000010000000011100001000000001000000100011000000000010000011000000000000000000001010000000000000010000000100000100001100000100000001000000001100110001100100001000000000100000010101011010100100000010101000000000000001100000010000100110000001011000100100010000000010000101100010010000010100000100001100001010010010000010100010000000000100000110001000010010010000000100010100011000000000010000110000001100100001000110000111000000110001001010000000001000000001000010000010001101001011100100011010000010000001011100001011000001100000100000001110000000000000000100010100000100000010100101100011001001010000000101110000000100110100000000000000010000000001000100000100010100010100100100100000110010001101111010001100100000000001000100101000001000110000000010000101001001100011001100000000010001001110001010100010110011000010001000000101010000110000000101000000001010000011111100000100000011001010001100000001001000101100010000101100001000000000011000000001000100000011000010000000100000000000000000010100100110000000100011000001010001101001010100100010000101100000000100101000000000100101001000000010000101000101010000000000001000000001000000000000101010100000000011100010000001001000010000000101100100010011010001000000010000101100101001100000000001010000001000011001100000110101010000100011010101000000010101100011000000001000101101000000001111000000000001000011100100000000001000000010101000000000110000001000100000000100000100110000000100000110001101000000110011001001001110000001000011000000000110100000010011000010010010000110100000000000000000010000100000100100001100101000001010010000000001000111000000010010000100000110000001010011000100000000100001001001000100000011010000000000000000111100001010100101000000000000011110100001011000001000101000001010011010000000100010110100000010000011000101100001100110100110001000110010000100001000000001000110101100000101110001100010000001100000000100010000000001000000000011000001100000011001101010100000011010001001000000100001000001001101100000000001001000010000100000010000000011100000000000011100000100000000000000010000000010000000000011000000100010110000100000111010000100110100000000000001000000011000001100010111000100001001000000000010101100000011001001000000110010110000010010100001000100000001100000000011000000000000000110000100000101101010111000101000000101001100000000011000110100010001000000100000011001001001001110010010001100001010100011000011001000011000001000000000010000100000000100000000111000100010100010001100100000000010010000010000111000000100101000101000000011001000000001001010000101110010000000001001001100100000000000001011010000000011000000100010001000000000011000100100100000110000010000100000100010100000001000001010001010000000010010000000000001000010110000011000011000010110010100001001001111000111000000101010011100000011100111001101000000000100000001000100000000000000000010011001001011100000001001000101000010010000000000000000101001001000000000010010010010001001101001100110100101000000100010001101101100000100001000000000100100000001000000000010000000000001000000100001000000000101000000000100011001100010001100110010100100010100000001011000000000000000001000100000010000000010001100010001000000001011000000011110000101000000101100000000110000000100001110110000100010010011101010000000000010100100011010101010001000100001001100000100010000101000111011000000010101001000100011001010000000000000001000010000000011000100001001100010000000010010000010000000000001000001011000001000100001010001011000000000100000000000100010010101010000000000010000001000010000001010100000000000000000010000011110000000100000110010000000100000101001010001000010000100101010000000010000001010110000100001000101101001011010001011000000101100000000110000000011000000000010000000100000000000110000001010101000000000000110000001010100000000010000000100001100010100000100010100000000000011100001000000010000000000001011010100000111000010000011010001001001010011010001010000101001001000000010001000000111010010100010000000010000000000000011011100000110000000000101000000000100100011101101000000000000101011100000010001101111000010100010110000000100010000010001110110001101010000100000001000000100000000010100000100000001100000000011001110000010110001101101101011100000000001000000100001001000010011100000000001000001001110010000010000000000000001001000000010000010000001000000000001000000100011000010000110010110000011000010000001110010010100010000001100000000001010010000001000000000100000001000000010000000000011000000000000000100000001000000100100100000100010000000000100000000000000101100000001100000000100011000011000000010001001100000100001010100010010000000010100000000110100110000010010010001110000001000110000010010111110000011000000000000111000010000111100000011000000101010000000010000110000000000000111100000001010100010100001000000000100000001000011100011000000000100100011100000110101100100011001100010000011010000111010001010000010100100100000000000000000000000100000001101111000000110000010110001001000110000010101110000000000000100000000001100000000010000010010000000110110110001110000100100000100010000001000001000010000000100010010000000001000100100000001100001000100000000000010001001100000010100010110000000000001100100101010101110010111011000010000000000011000000000011100010000001101000001000110000000001000000000000000000100000101101100000000000100001010000010010000001000000000111000000100100110010000001100000001000010001000001000000000100000000101011011000001110000100000011000000001000000010010000100000000100100101000100010010000011010000001010010000000110000000000000000000101010000100100010000000000000001100001010000001001101000011100000001001000101000010010000000100010000101100000000010010000001000000111000000000010011000000100000000111001010101100000000101011000000001001010001010100010000010000000000010000011010000011000000000010011100001010000000000100010100000000100010000110001100000000000000101010000110010000101111000000111001000001110000000011000000000010000000100001000001010000100000101101000000000010100001100000101000000000101000001000100000111100000000010000100001000100000001011000101001100000000000010110001110001010100101000011000100100000000011000001100001101001001011000000100100001000000100011001000000010010000010100001000100010000011010001100001001000010110000100110010110000100001000010000000100000000000001000001000111000000111010000010000001010111001100000010110000110100001000010010010001000000100010000010100000100101001000100110101000001000100000100000000000101100000000100000000000010000001001000001010100001000000000000001000000011100000011000000000000100010000000000010000110011000010100110000100000001000001001010000010000000000001100010001000000000100000000010001111001000000010000011000000000001000000010001110100010000000000000000010100100000100000000001100100000000001001110010100010000000100000000001010000011001000001000000001000010001000110010000011001001100101010000001001000000000001000000101010000000010100000010001000000000010001111000100000001100000101000000110001100000000000111010000000100110100100001100001011000010001000001001100000000000001101010000010000001000100100001011000000000000000010000000001000001100000000111000010001011001000100000000000000010010010001001000100001011000100000000001010000000000000011010001000010101000000001001010101011110000000000001010000010000000011100000000000110010010000100000001011010000010110100000001100000100000001000000001000001000001100100000000000000010001010101001100000000010101000000000000000100000000000000001000110100000001000010000100000001010000001100000101001001000000001010000000010000000000001100000011000000001001001000001011100010000000000000000110110001000100000000010000000000110001000110001010001100100101010010000001010000101000011001101010001000000000100000000100010001111000110000001100110100010000000000000000000110100100001000000000001100011000001000010000100110001000000000000001100000000011110100010010011001100000001100110010001000110110000000010000000001100000000110001000100100011010000011000001000101100010110000100000001000010010000000010101000000000001100101000110000100000001000111000000",
	"1111010000010010000100000000100000010100100001011100011000010101100111100001000010000001010000100100101110001000000100000001001111000011111000111000011010010011100110000100100011011001001001001000000110000001000000000000100101010000001000000001011000001010000100000001001000000100101000101000111000001111001001000100010000000000001110000000001100001001000000110000011110110000110000001000001000001000010000011101000110110101110010001000000001000101000100001110010001001000001001000000000000100101101001101000000000001000010000100111000000001000000000100000000000000000001101000001000010001010110000001000010000110001001110000000100000010001000001000001000010011010100000110010000000001001101001100100001010001000010000000011000100000010001001000001100000001000110011000100000101100010001010000001000111001101001000111101000011011100001110010101001000001000000010000010000000000010100001000000001000000010000000000001001000100100100100110001010000010010100100100101110110100000100111101001011000110101000000001001000000100101001001101001011011011110000001100000101000011000101001010000101100011101010000110010001001000110010100010000001001011000000101000000000000000000010100000110000000000001100110100100000010100101001011001000110100001000010000100001010000000000000000010001100100111001111011001000000101110000000010001010000100000001000101000000010000011010010001001001000001010001000100100000000100000100000000010010110110100010001010001010000001000000010000001001000000000100000000100000100000011000100011100000000010100000100000001010110000000000111100101000110010000000001010110000010010001000100010100011110111010000100100100010001100001000010000010000100000000000100000100000000000110000000000100010100101001110101000100100000100000001100100000000000001001000000001001010001001001010000000000001010100100001001010000100000101000000110101000100000001001100001011100110000000010000011100010000001000110010001010000110001000001000000000000000011010000000010000011000000000000000101000000001000000000010001000000000100000101001100101010000000001000110010100110000100000100000000000001011010100100000011001000000100000001110000011000100110000001010100101100010101000000100101000011010000000100000000101100001010010010000000000010100000000000000101000000011000000000000100010100001010010001010000010100010010010001000010000111110000010000101000010010001000100001010010000010000101111011100100001110001010000011001010000000001100000001000000001100000000000000000000110110000100000111101001100010000001010000000001000000000000001100000100000100001100000001000100000101010100001000000000100000011010000001110010001101100000000001001010101001000000101000000010000101101000100010001001000000010001001100000000001010100001000000000100000001000000101001010000000001010010000011011000000100000001000010001100100001001000100000010000001010000000000100011000000001000100000010001000001000000000000000000011000100100101000100100011000001000001100001010100100010000101100000100100001001000000110101010000000010001001000101010000100000001000000001001000000000101000100001100010000010000001001000000000000111101100010011000001000000110000101000001101101101000001000000000100111001000101100111011000101110010001001000001001101110000011001001101101100000000111000000000101000010100010000000001000100000101000001000001000001000100000000000000100000000001100001110001101000010100010000000001100000000000001010010100100010000000000000010100000100110100000000000000000000000111000100001001001000000101001001010001101000001000000010010100100001100000011000010100100000000000000001001000100100011010000000100000000111100001010000001000000100000001000100001011000001000101000011101011010110000100010000000000000000001001101100001100100001110001010101000000101101001000001000110100000000000110001101000000001000101000000010000010000100000000010000001010100011000111010000001011010001101000000100101000000000101100001011000001000010010100001010000010101000000000000011000000100000000010000010000001011000010000010100000000010110010000100111000001000110100000000000001000000001000000000010000001000001100000000000010101000001111001000000000110010000000010010010001000100000001100010000010000000000001000100010001000011001000101100101000000001000100000010011000111100000001010000000000011000001101000010010010000100001001000010000010010000011000000010000000110000100101000000000000110000101011000010001000000000000010011000001000111000000100010000100000000010011000000000001010010101110000000000001001001110100010000010000000110000000110000100101010100000010010001000100100000010000000011000100001100010001000000000010011101010001000010000000000100001000110110000010000001100010010010100000001101110000010000101100010011011000001101111101100010000000100100011010000000000001000000010001000011001100011001001000000000010010001000000100100100000001000010000010100100010011001100000100110100000010000001010001001111100000101001100100100110000000001000000000000000000010001000000111011000010101101001000100100101100100010001110100111100010011100000011001001000000010000011001100000011000000010001100010001000000000001000100011100000101000000011100001000010000000100000100010101100010110001101000000001000010000100101001000000001000100001001010000001000110101010110011001101010011000100000011010010100000000000011000010000000010110100010011000010100000001010000010000001000011000001001000000100001000010001011000010000011001000010100010100100001010100100000000100001010000000000010100000000000000000010011100000000101100010000000000101000001000010001000000000000100000100000010000001010110100110000010100101000011010001010000000000100010100000000000001000000000010000100100000110000100000010000101000000010000010000001110010001000010100000101000000000101100110010100000000101001001101010000010000000000000100000001000000000010101011010011001101010011010001100000101011001000000110111000000110010110100000000000000010100010000010011100101110111000000110000000000000000011001100000000001000011011101000010001001010100000100000110000000000000000010000110000101101010000000000000000000000100010010100000110100101101100000000101110000001010000101100001001000000000100110000100001000011000010101000001000100100011110011000001000000010001001000000100010000010001001000001100000000001100001100010000110010111000011000010010001110000000000000111001110010000001100010010001000000001100000000000000011000000000010000000000000010000000001001001100100100000000010001000000100010000000000100100000011000000000100011010001000000000000001100100100000010100110000000000110000010000100100110000010010010001110000000100100000010010010110000011000100001010011000010100010000000011000100101110000000010000010000000010000111110000000110100011101011000000000100000001000101001001010001000000100011000000000001100101011001001010000010010001011010001000101100000100101100000001000000000000100000001101100000000110000010100000001000110100000001001001000000000101000000001000110000010000011010000000110100110001010001100100000000110000001100000100010000000001101000000001001000100100000011000001100001110000000010000001010000000000010011010000000000100010001000101110000101010001010000000000001000100010011100000000001001000000010010011000001000100000011000100100000110110100000000010100000010000011011010001010001000011100110100000010010100000001010000100011001000001000100000101010100001100010000000110000100000001000000001000100000001000110010000000100101000001010010000111000000000010000000000111000000000101000100011010000000000000000100000000001100001010000011100111000011100000100001010101010010000100000100110000000000100000010010000001000100111000000000001010000000100000100110000010001100000000100011010000000101000001110100010001010000000001010001110110001101000100000100011000001010000000000100000100001000001010000110000000000000001000100010000010000100001100000000010001000001111000100000000000000010000000100001000001000000100000101001000000100001100001100000111000000000001000001010000000010100000000010000100000010110000001001100100001000000000001010110000101000010100000001000010000000000000101000000100000101001011000000010100001101000000000001100000000010010000010100000000101000010100000011001001000010110001000000010010010000101001100010010000100001000000001001001000111000000111010100100001001000110000100100000010100100000001000000010010011000000101010000110100000100000011100010000100000010000100000100001100000111100000000000000011001100000001001000001011100010000100000000000101000011100000011000000000000110011000100000010000110011000000100010101010010001000001001010000010100000000000100000001000100100100000000010001011000000100010000001000000100100000000000001100001000100000000110000000000100000100010000011100110000000000011000010010010000000100000000001010001011001001001000011100001011001000110010001010001001000001000000001011000000000001001000101100000000010100000001011000000010010001001000100000001100000111101000000001101000001000101000100000101011100100010100001001000000001000001111010000000001001110010000000101000000100000001111000000000010000010000000100100001100101000110000000000011001010000000000100000010010010000001110101101010000000000000001110000110000100011010000010011001001000001000100101100010000010000000010000010000000010001000000000110000010010100000111001011100011000100000000000100100101101000000001101001000001100100100000101000000001010101001000000000110100000000000000000000000000000010000010010001000011000010010100000000000001001000100100001001000000100011000000010000000000001000001010000000001010000000000001100010000000001100001100010001000101100000110001001000110000000111000010101100000101000010010100010000101100010000100001001010010010000001100100010001011000010001110000010100010000000000000000000100100110001010010001000100011000001000010000101110101000000000010000100000000001010100100000010011000000001110110000101000110010100010010000001000100010000100000001100000011010000001001000100111100010110000000100001001010000000100010100000001000001011100100101000100000011101000000000",
	"0001000001010100000000000100100000000111000101010100010000010101100000100000000010001000010001000000110000011000000000000001010001000111110101111010011000010001000010000100100010011101010001000010000100000001000000001000000100010010000000100000101000100010010100000001100000001101000000100011011000011101001001000110010000001000001100000011001100001001000000100000011110010000100000000000000000000100000000010010000010000110010010101101001100010001000100101000010001001000100000100101000100100001101001101000000000000000010000001010000000100001011100100000001000010000000100000000000100000010010100101100010000010001000110001000000000010010011101000001000010001111111000110110000000000000101100000100000000000100000000001011001100000000011001000010000000100000101000000000110100101000011010000001100110000000000000111101100111001100011100010100000010000011000011000000100100000010011001000100100010000011010000000001001000110100100010000001010110110000000000000101010010100001100001000010011000001101100001001101111000110000001000110000001001010100100001000000001000011000111110010000100000000100010010110000000101010010000100000000011000101000010100000000000000000000010101010111000001100001000000110101010000000001111110100000110000001010010000100000010000100000000000000101000110011101011011001000000100110000000011010111010000000111000101010000000001011010000001001001000001000000000100100000001000000100000000011000100000100010001000001000100001000110011000111001000000010000000001000000000000010100000010001000010010100100100000001000100000000000101100110000110010000000001010010010010010001010100000100101010010010001001011100011001000010000100000000001100000000010110000101010000000010000000000010010000101000010010001001000000100000001110000000000010000111000000000011010000001001010000000000000000010100111001000010100101100000010110101001001110001000000001001100110010000011001011100110010000000100000011000000100100100001000001000000000010000000000010011010000000001000000001000010001000000000010001000000101100000010001100011001000000001110100011100000010100001000100000010000000010000100000000101000000000000000100000010000100100000001011100000000100000000001100000000001000010010100010101001100000010000001000010001000000010100100000010100000010000000100000100010000101000010001011010110000011110000001000010001100000000011001000000001000100000100000001010010010001001111110001000000110001000000001000100001100001100000000000000000110000000000000000000100010000100000011001001100010000000100000000101110000000000011000000100000101011100000000000101110000010100000000000101100010001010001000011010001101000010000100000110001000001000000000100000000101110000100000001111000000000001001110000010101010101000000000000100000111010000100000110101000000010011000110011000000011001000000000000100110001000000100000001000000101000000000100011000000001000001100011001000001000101001000000000001000000001111001100110000000001010000100000110100100010000001100100001110101001000001110101010000000010001001000001000100000010000000000000000000001000111001100000000010000010000001000010000000000111101000010000000001000000010000100000001001100100000000010001000000010101100100000100000000000011010001001000010000100100110010101110100100000000100111000000000101000010100010100000001001000000011000101000000000000000100000000100010010000010001010001101001101000000100010000001001110001000000000010000100100010010010011000010100000100010100000000000100000110001011000100001011000100000101001001010000001000010000001010010000100000100000001010010000000000010100000000001010000000011010000000000000000110000000010000100000000100000001010000011000011000000111000001101011010100010100010010000000010000000011000110001100100101000011010101000000000001010010001000010100100000001110000100000000000000100000100010000000000000000000010000001000000000000001011100000110000001001000000100101000001000011000000011001001000010010000000010000000110000100000000011001001000000000000000000000001010100000010010000000000010100001000000100000000100100100010110000001000000001000001000010101010000001100010000000010101000000001001001000001110010110010010000110001000000000101000000000001000000000000000101010000001100101000101100101000000111000100000010011000101110000010000000000000001100001101000110000010001100000111100010001010001000011000000000000000100000100110000000000000010000001011010010001000000000000000011000011000100010000100011000101000001111011000000001011010000101100010001000001000101110100001000010000011110000000010000100000110001000000000000000001110100000010000010000100001000000101000000000101011101110000000010110000000000000000100110000010001001100011110010100000001000000010010000100001010000011100011100011101001000000000100100010000001000001000000000000001001010111110001001001100001000010010100000000000010101100001000010000000100000010001001100011100010100100000000001010001011111100000101000000100100000000000001000000000000000000000000000000111001000000000101010000101000010100000011001110100111100100010000000010001000000010010000010000110000011001000010000100110000100001000011000000100010001001000100111100010001010000000100000110000100000010000000001010010001100000000000000010000000000000100001011000000100110100101010101001000111110101001000100011000000000001000010010000010010000000000100001000100010000000001010000010000001000011000000010000001000001000010000011000010100000001000010100010000100011000000100010000101000100000000000100100000000010000000000000110100000100000000010000000101000100000010001100010000000101010010000001100001010001001000001001100101000001110000000000000001100011100000000000101000000000010010000101000010000000000000110101000110010000000000001010000001000000000100100000100000101101010100110001000001001100010000000000000000000000111000001000110000010111011000011001101010011010010010001101010110010000110100010000101000010000110110000010010110010000001010100101110010000010001000000000000000110001100000000001000110100101100000001000101100000001000010001000000000000000001100101101001010010000000001000000000101001100100000010000100101100000011111110000000010001100101000001001000000101100000000001000000000011001010000000000100011010010000011000000010100000001000100010001110000000000100000001000000100111100010000000010110000011000000010001110000010010000111001010100000001100010110011000000000100000001010000010000000011001000000100110011100000000001000100100000000100010000000000100010000000000001110000010100000000100011001010000000010001000100001000010000100100010000010000000010000110000010010010000010001110000001000110000100010100110000011000000001110001000000000001000000010000000000110000000010000110000000010000111100000011010100010100011000000000100000010001010100101010000000100100011100000100001100001010001001100000010010001101010001001000110001100101101000001100000000000100000001101100000000111000010000000001000110100010101000001000000000101000000000100100000000000010010000000110000010001010000000100000110010000011100001000010000010110010010001000011100001100000001110001000000010000000000100000010000010000000011011000010001101100000000101110010001011001000000000000011000110010110001010001011100000101000100010000001000000000011000100000000100100100010000000000000000000011101000001010001000111100110000001100000000000000001000110111001000001000100000101011011100010000000000000100100100010100010001000000000010010000000000100100101100111000010000011000000101000000000000111000000001100000000101010000000000000000000000000001110001010000010011010010011101000000000010101010010010100000000100100101110100000010000000000000000111010001000001011001000000000000100000010101000000000101011010100001001010000011100010000010000000000010001001110100001001100000110010100000010101000100100110000001100101010000110001000010000100000100011000110000010001100010000101001000101110000100010000010000010100000000000000001000110100000001101000000110000000000100000101000000000000000001010100000010100000000010100100000010100010001000000100011000000000001000100001111011010110000000000010000000010000001000101100000111001010111000100100001110000000001010100000000000000000010100000000101010000000010010101000001010010111010100010110100000101001100011000000010011000000000000000010111001010111010100110001000000111001000100000110000000000001000000000010001001000001010000010000000101100011110011000101000010000000010100011000000101100000110100000010000000000001001000001011100001000100000001001000101001000001011000010000000000111000000100010010110010000000100110101100010100000000101010100000100100000001000010001000000000000000000010001110000000101110000000101000000001000000000011111001000100000010110010010000010010100000000010100100100000101011111011000010000001101000000000110001011000000111100010001000111001100110010100001011000000100000000000000000000000001000000101010000000010000000000001000010011010101101101100010000100100111011100100001101010001000110010000000101000100101011100001010100000001000001111100000000001000010000000010000000000100100000111010000000010010010000010001000101000001000101000100011011000110100000000100000010010000001001011011001011000000000001001010000100000110000010000010011101001000001101000101100100000000000000000000010100010010001000100100010010010000101000000010000000001000100001001000000100001000000000001000000000001110001100010000010000000010100001000000000110100000000000000000100000000000011000010000101000010000100010000000001010001000100000111001011000000100001000010110000101000000110000000000000001001110000001011110010000010000101000000010000000000000000000000000000010001010010001000101100000100000010010001010000000110011000000001000000110000101000000000000001111100010001111000010101001000000011000001100100101110001110000001001100011000001001000000001110101000000000010000100000001011110101110011011000000000001110110001001000010010000001001000000000100110100100000001110100110000000001000000000000001000100000100100000001010010000000000011000101100001111101000101000000000010001001010000"
	); --six test class HVs, one for each vowel
  	variable test : testarray := ("1101010000010010001100000100100011111111110001011000011000000100100010000000001000000100010101110100100010011001001100000010000010100111011000011010001010010010000010000101000001011000001010000011010000000001001000001000100001010100101000000111001100101000000000000001000000000000001000100001111000110110101001000110010000000000001111100011000100001000000010100000001100010000110000001010001000000000000100001001000011000000001000001000101010010111010001001100010001001000011001100001000100100100101001000000000000001000001010100101000000111110111000000100101000010000001001000001000110001000110100000100000000000000000100011000100000010000001100000000000010000000100000000000000000001001111111000100001110101000010000000001000000000000010000001011110010101000110010000100010001110010001000000001000010010001001110101100000001001101000101011101001110100011000011100010000100000000010001100100101001100010000000000101001100100000000000001000000000101010101000000100110000101000000001100011011010001101100001000101100000100000001000100001011111111100100010000010100101001000101101010000100100011101010000010010001100000010010100010000001101011000010000000000101000100000000100000001000000000101101100100101110110000101101111101010010100000000010000100010011000101000000000010001000110111000110001000100010000010010000010011110010000101001000000010000000000000010010001000001000000010001000000100000000100000000100000001110100100100000000010001000010000000000011100011001000001000000000000110100100000001000100000001000010010100000000000000010100110000000111100101000101010000000001000110000000010001000100000100001010110010001000110100001011100011010100000011001000000000001110000000010100000010100100000100000100000000000011000000000000000000011000100000000000011101001000000001000001001001000001000000000010100000011011010000101001001000010100101000001100101001100000011000111001000010101100100010010101000010010010011000110001101000010101000000100100000000000011011011000000000000000001000000001000000000010011000100000100001111001100000011010010001100000000000100001100000100100010010110001000000100100000101000000000000001000000001000100110000001000000100100110101011000010001100010010011010100000001100100001110010010000010000010100000100100000111101011000010010000000010010100111000000000010000110100000100100001000010000111100000001001001010010000001000000001000010010010001101111001100100001011001010000000011100001001000000000001101000001010000000100000100100000101000100000010000101000011000001110000000100010001010100110100000000000100010000000001000100000111001100011000000100110001010000101000011010001000100000000001001110101001001000110000110000000001000001000011001000000010010000001010100010100010100000000110001000000111110000100001100101000001011000000010110000000100001010111000000100010010001000101100010000101010001100000100100000110001000100100011000010001000101000001000000011010100101110000000100010000000010000100001010100100010010101100000110100101000000100100000000000000010000101100000010100001100011000000000000000000000111000000001000011100100000000000010000000000001100100010010010010000000000000101100101000001010000001000011000000110000100000110110000000001100000100000000001000111110000000000100100101100000000111000000000001001010000010100000100001100000101000101100101000001000100000000000000010000000000100000110001110010010100011001000001100001001000011010000000010010000000010000000011010000000110000010000100000010000000000100101011000101000101011001010100001000111010000010010000110001010000010010001100100000000100001000001000100100011011000000100000000010000001010000101000000000000011110110000011011011000111100011000011000110010101010110100000010000010010101100000100000001110010000110010000100101010000001000101010100000100100001101010000000010000000000110101000001000000000011001011110100011000110000100000111000001011100000100000000001000110100000010001001000000000100001010010000001100000000000010100000100000000000000010000000010000010010011000000100010110010100000000000000100110100000010000001000000011000100000010000011000001001000000000011101000000101000001000000100010100010010010000000000100001101100110000010000000000000000011010001000111001010110000001000000101001100000010011000011100000000000000100000011101000101001010011010000000000011100001100010111000001000001000000000000000101000000100000000101100100000100010000101100000001010011010000000111000001110110000101001000001000000000011001110000001110000000000000001001100000000010000001010000000000111000000100010000000000010000000100000000000110000001000100000100010100000001000010010001000000000010010000100100010000010010000001000010000100110010100001001111101000111000100101000011100110001000010100000011000000000100000000100000000001000001000011001001111100010011001000000000000000010000010100100000101001000000010000010100010001101100000100000000001010000100010001001101000010100001010000000110100000000100100000010000000000101000000100000000000101000001000100100011001100000101000110100100110000100000010000001100010000000000000100000010000000010001000010001000011001001001000011110001100000000011100010001110000001101000100110100100010110110100010000001000010100100010010011000000000000001001000000100011000001000111011000100010010000100010010000010000100000000001000000000000010000010001101000000100000011010000000010001000010000101011000000010100011011001010000000000001000000000100010110101000001000000010001001001010000000100110000000000010100010010011000100000101100110000100000101000001001000000000010000000100000100000011100001000000100100001011100001001011100000010000000101100010000110000000010000000010010000000100000010000110000011100101000100010010110010000010110000000011000000101001100000000100101010010000000000011100001000100010000000000001111010000000110000000000011000001001101010001010001000001001011100000000110001000000111000010110000000000010010110000000011010000000010101100000011000000000100100110000001001000100000101011101000010000101111000010000000110001000100000000010001110010011101100010100001100000000000100000110100010110000001100100000011011000000011110000100101111110101001000100100000000001001001010010100010001001000000011000101001011000001001000001000000100000001110010001000001100000000001100001100010001000010111000011000011010101010010010000010110000100000000001010010000001100000001100000001011000010000000011011000000000000000000000001000001001100000001100010001000010110000000000100000000000000100000000100001000010000000011001001100101000000010100010000001010010000000010110100110000010010000001110000000000100010000011110000000000001100001100011000011100111000000010000100101010000000000010010000000010000111010000001110000110100001000010000101000001000111101000000000000000100011001000010101100111011000101110000010010000110010001000001000100100001100000000000000000000100100001100010000000010000010110011000000010110000100111000000000000100000010001100010000010001011010000000110110000001000000000101000000010000001100001100000000010001000010000000001000101100000000000001100100100000000000101000100000000100010111000000000000100110000010101010111111011101010100000001000000000000000100010101010001000001010010010000001000100000010000000100000011101100000000110100000010000010000000001000001000011000000101101110010000000101010001010010000000001000000000101000100100000001000010010000100000000100010000000100010010000110000000000000101000101010110000111000000000010010000000100000000001001000000001010000100100010001100000000011000001000000010100111010011101000100001010001000000000001100000111100100110000000010010000001000100000000000000000011000000000000000111001010000100000000101010100110001011000000110000001000100000010010000001001010001000000000000010000001001010111000001000100000000000001000000010001000000000000000000000000010110110101011000000111001000000111000100001000010000000000000000001000011011000100000100101010000110011100001100010010100000000101000001000010000100000000000010100100000000000010001011010101001100100000000000100000010010110100101000000000100000000001010100011100101100010001011000000100100111000000100011001000000010010000010100000000101010000100010111101000000000010000100000010010110000100001100010010000000000010000001000011010001001000100000000110001001010111001000000010000000110100001001000010010011001000000010000010000000100001010010100110001000001000100100100000000000101100000000001010100000110000101000000000011100011000000000000001001000010100000010000010000010100011000000100000000000010010010000100101101000001000001001010000010100000000011100011000000100100110010000000001101001000000010000011000000100000000000000001110110010000000000110000001000000000000010000001100000000000000001110000110000100001101000000101010000001001001001100000001000011001100100010101010000011000001010000000010000000000010100000101110000000000100000000011000000000000001001100100000000110000111010001100000001010001000100100100100101110100100011000000011000010001000001101110100010000001000000000100000000000000100001010000000000000000010000000001000001100101000101000000101011000100100000100000000000010010000000100000000010000100000000001110000000001010011010001010001100010000000001000001011110001000000000000000110000000010110100100000110010000000001000100011010000011100100000000110100100110000000000000001011000001110101000000001000010001010100000100001000010100000000100000000000000000000000001001110100000001000010000000010001010001001000000100101001000000001000000000000000101000001000000011000000100011001000001011010000000000001100001111010001000100000000010000000000111001000110001000001100100100010010000100010000100000010000100011001010000010100000100000000001010000010000001100010100011000000000000000000100000010000100010001001100010000000000010000001010001000000000000010000000001111100001000011111000000010000100110110000000110101000010010100000001100000000111101000100100000000000011001001100101100010010000000000101001010000000000010101000001000001100101100110000100000001000000110010",
	"0100010000000010101100000100100010001101000100011100001000000000000001100000100000001101000101000100100100010001000100000010011100110011101001011010001000010001000110001000000000011001010000001000010100000001000010001000000100010100100001000101011100001010000000000000100000000100000000100011110101010101101101000000010000001100001110100011000001000000000000010000011010010000010001000010001000000110000100110010000010100101000100000001101100000110011101100100100001000000001001101000001110000000100001001000000000000000000000000110000000101110001000000100100100001001001001000001000110001010100000000000000100000001001100010000100000010011000101010001000010000100011000010110000000000001101001100100000110001000000001001001000000000010011100001011110010000000100001000100110101010010000000000010001111010101001000100100100111010000010011000001001100001001000001000000000000010010011000100100101000100011010000011000000000101001000000100000001000101010001000100101110010000100000101000011011010011101000000000100111000010100001001010001000011001100000001100000100001001001001000010000000000010100001000111000000001000100010000010000001001010001001110000000100000000000000100000011000011100100101110100110110010100100101110000010100000001010010000000011010000001000000000010010111000001100000110001000100101000010000001010011000000001000000100010000000000001010000000001000000001000001000001100000001100010000100000010000010110100010000010000010000000000000010101000000000000000100000000100100000000010000110001101000000000100100100000000010100010001000111100011000010000000010100000110010010000011000000100000010010000010000001101000011011000000000110000010000000000010011110100101000100000000000000000110010100000001100011001100000100100000000100100000000010001101001000000010010010000000000000000000000000100100010011000011000100101000000010000001101100101000100011000100010001000001101010000001010001000110010011011000101000001000010000000000100111010000000000100011000000011000000100001010000000000000000011000100101001101010001000101011010010001100110000000100000100000100000010000010001010100000100000001000000000010101010000001000100000000011011100001000110001001011000101000010000001011100000100001000001001000011000001000010000010000000000110000000000000010100000000000100100010000001011010010100011010010000000010000100010000110001100010010010101010000000000010010010100000110100101000010101001000000110001000001010001001110000001000000010000001000000000000000100010110000101100000000001000000100000000101000001011000110000000000000000011000000001000001000010000000001100000001000110000010101101101000001100100000000001000100100000001000110000010010000001000000000011000110000010010000000010001010000000000011000110011001000101100000110001000010000000001011000000011000000011000010010000000100010001000000100100011000001111001100000000110000100001000100100001001000101000000001000000000000010100100000000000010001010100000000100000000000100010010000000100110110100001000000010001111000000100000101000010100000000000001000100000000000000000011011101100100001000010000000000010000000000000100100010001000100000000000000000000101101101001000001000010001100110100100001100100011000100111000000001000011101100010100001101001101001000000101101000000001001000010000000000000000001000010010010001000101000001000000000100100000010000010001010000100000010000000000000000001000110001010000011000000000010100010000010000010100010100100010010010000100000000000000000100100011001000000000001001000000001000100010101001010000100000010000100010111000000000010100001001000111000000011001000000100000000010100001000100000100100000000000000010010001010010000000000010000010010110010100010110100101000000000001001010001100110001110000010011011000100101011000001000000110100000101000000101010000001000001000000100000000001000000000000000000110100010001101000000000010000001110010001000100000001000011100001001000000000000011100001010000010110100100100000000001001000000001000000010000000001101000000001100000000010110010100000101010001100110100010000000010000000011000001100010000001101000001000001000000101000001101000000000000100010110010000000010001000100000100000110000010100000000000000111010000000010000000011000100000000001001000000010001000101100000010000000010000000101001000000010010010001000001000100010101000000000011000001010000100100000100000000000100001011000000000110010100100100001000010001010011000000000001000100000001001001110000000000001010100010101100010001000001000101010000010000000001010000000000000000100000100001000000000110000000000100000000000000100100000000010001000001000100001001100000000000010000100000001000010010000001000001100010100010100100000000100000100000001100000010000110001000111011110001000000000100001000001000011000000001000101001001111110010000001100101100010010010000000000100111100000000000000000110000010010001000010100110100000010000101000000100011000000100001110000100100100000000000000000010000000000100000100101011000000001101010000000100111100000010101010100011100010001100000010010001100010000000010001000000011001010010000100110000100001001001001100000111101101001100011000011000100010000001011100010100100000010011100010010001100000000100011000100011000000000000100110010101101010101010110000000000010101100000000001011000000001000000000001010010000001000110000001000010100000011010000010010001000001000101000000000110100011000001011100010001110001000010100100001100011010000100010000100001110110001110110000000000001100010010011010110100001100100010100000100000000000000001000010000000000001100000001000000010000001100001001110001001010110001001000000100100010101110000000011010000010000000000001000100000000000001100101000000010000110010001000000000000010100000000011100010000001001000100001001100010100011010000000000000001000001000101011111000010011010000011000101000010000001110001001000101000000000110010000000000110000100100000010000110000000010011100001010111000000001000000000000100101100001000000000100111101001001100000000000000010000010000001000100000000101001100011000001010000000001000000100000001000000100000100100101000000000000000000000000000001100000100101100000000001000000000001001001000010101000001000001101000010110010010000001001111000000000101000001110010000000100100000000001100011100010001010010111000001000001010100010010000101000000000010110000001100000100011100000000001000001011000001000000011011000000000110010001000001001001000000000001000010001000010100000010000100100000000011100000000000011000000000000000000001100101001010010100000010000010110000010000000010100010011110010000010000000000000010010000001010000010000100001110010000000100001000010000000100001110000000011000100000000000000000000000011100100111101001000000000000000001001011000111110000000101000001000000100000100001001001101000000011010001110000000001101000000000000101010000100000000000100100011100010100000001001000110001001000100011000001001001000000001101000110001100010000010000011000010000110110011000100000100000000000111000011000001100010001010100001010000000011100000000000010100000000101010010000010001001000000010000000010001000010001101100101010100000001111000000000101000001010000110010100101000101001001000101011010000000000000000001001000101110000001011100010000010100000010000000110000000000000000111000100000000100000100001001011001000001000000000000000000100011010000101001000010000001100000011100000100000100010001000010000000100001100100010100000010100010000110000010000100011000000000000010100101010000100100010000000000000000110000000000010101101010011100000001000000101010000000001100000001100000000100000010010000001001100101000000000011001000000000000000111000010100000001000100011110000000110000000001111110000010000000000010001110100001110100100000110010000000000000000101000000000001000110010000100000001001000101000100000000010010010110011010000100000000100111000100011000010000000000000100001000010000010100000001001010000100000100000100000111100100100101100001000100000110000000000000100100000010000000000101110101000000000000000000010001001001000010001000101000100100000001110100010000000010011000001000100000100000000000100001101000000000000010000000000000001010000110000011101001000001010011000000000000100010100000000011010000110010000000001000011000001000010101010100100001001000111000001000000100100010100001000000010010000001001100010000000100001000101000010001010001100011000100100000001101000011100000110100010000001000000001001000000000100011100110000001001101100001000101011000010000000100100000000000000010110000000000100000101000000101000110100000100010100100000001000001001000100000110010000010000000000000101010000001001000000001000000000110101011010000000010110010001100011011100010000000100110100000101000100000010010000001100000000000000001010011001111000011000000000010000100010100000010000000000010100011011000000000100111000100100000110001000000011001000010011010101010001000010001100100000110001000001100010101000000110100000000100000000000000000001000000000000001001010000001001000101011000110101000000001100000100010000010011011000000010100000000100000010011010000000011000110000010100100010010010000001001010000001011000000000001101000000100001000000001001000000101010000001100110001100100001000000001010000000100010011101000100000000000010010100000100000000000011100000000000100100000110000000000001101010000001000101000010100010010000010001000000000000000101000000000000001001000000100000001000000110100001000010000100000000010111000101000001001011000000101001000011110000000001000100001001000000000000011001001010110010000000001101001110000000000101000010110000000100010001000111001000111000101000010001010000101000001010000001100011001000000000101000100100011001101101101000001100100101101000000001000001100110000100001010010001000000011000000000010000100010101000000000000000000000000110000000100011111101000010001100110100100000110110100010001110000001010000100000101001100000110010000010001001000010001101000000000000100001000010100001010101000101010001110100000011000000000100101010100100",
	"1010000000000000101000010000000010011010110100001100001000000001000011000001000010000001000001110000001110001001001100000000001100000011101100011010010010010010100010011101100001000001001011001011010010000000001100000000000101010000001001100000011000101000000000000001100000001100001000101000100101011001100100000000011000000000001010000010011100000001000010111000011000000000110000011010000000000000001000101101000111110001101100001000000000001000011101101010010001000000100000001001001000100000100001100000000000000000011000100010000010011010010000000100100100011001001100000001000110001000010000001000010000110000001110101000000000000011010001010000000010000000100000010100000000001000010001100100000010001100010000000000001100000010001101001010110010000000010001000100010000110010000010000001001001010001001010011001000001011001011011011100000010000010000001100100100000000010111001000100100001000011010000000101000000110101000101110000010010000010100100000101010000101100000100101011000010101100000001001100000000110000000001011001011110010110000011100000000011011000110000000000111000010000000000000010001101010100000100000000001000110000011010000000100000000000010101010001000010000100101110110100010000100100100001100000000100000010010000000011001000000000010000000000100000010001011001000000010101100010000001001101010100001101000101010000010001001000000001000001000001110001000101100000001100110100101000000010100110100010000000001000000001000010010001010001000001010100000001110100100000010100100001000001010010000101100000000000100000001000110100111000100000000000100010010010010010001010000010000010110110000001000101000010000100010000110100000000000000010010100100101000100000110100101000110010000001001000010000000101000000000001110100000000010010101000000001000000000001000000000000000001010100000111010000000000000100000000110100001000000000001100010011100010001010010101110000001000001100110000000111000101111100000001100000000000000000000000001101011000000000000000000001000001000001000010011000000001100001011001100001011010010000000010011100010011000000100000100011011000000000100000011100000000000010101010000000000000000000000000110000100110101010011010001000010000011000100010000101100001011010001000100001010000000000000000100100011000000000000000000000000100000000000011000000100010000100001000000000101010000011000100000000010001000110000010000010011000100001000001000010111000000000100001110001110000101100001100000001100000001100000000000110100000001000111000100000010001001010000000101100001000000000100111100000101001100000000000101000100101100010100100000100000010000100001110010000101000010100101001010101000000000111000000010000001111000000010000011000010010001001000000010101010110011000110011000000100100000111000110001000101010010000000000000000011000001011000001100100010001000101000011000010000000100000100010000010001000100000011001000101000001001000000000001000100101010000110010011010100000101000100110100000010010001100100000010001000010101100110111000000110000100000111000100001010000000000001001000000000110011101010100001100000000001001000010000000000111100000000110110000000110000000000101101001011000000000000000100100000000101100001011000000100000100000000001000001001000000010010001001100000101001000000000001000001000110001000001000000000010000001001011000000000100000000001010000110010100000101101000000000010110011000000001100000010000011010000000000000000000010000000010000100010010110000100100000010000100000000000010101000000001010000010000100000010010101011010100000000100000011000100100000001000100000001001100100100011000000000000000000010100001010100001100100000000011000100011011001000000000100011000001010110000100000101000100000000000011101110000001000101000001010100000000100000001010000001100000000000100000101001000000001101101000100000001010001110000000010000001000000011001110010000001010000000001000001100000000001001110100001011000000100000011000001010010010000100000000000010101000100000001010000000100001001001010010010000000100110000011000100111000000000100100010100000001000010000000100100010100100101000001010100000010100000000110001001000001110010100000010000010001000010001000100000000001100000000001100110001100000100000000010110101000000100001100000000001000111000000011000000000000011100001001000000000000000000000001100001001010100000010000001010000100010001000011000000100001111100101011000000000001000000001000000010001000101000000110001010000001001010011000000010011010010101000000000001001001110100000011010000000000110000000100000100100000001000000010010000100000000100110000000100000001100010001000000000110010100010000000010000000000100001000100110000010000000100100100010000100000100100010011000100100010000011000010000010110110000000010100100010010000000010000000000010101001001101100001011000100100100010010101000010000000010101001000010000010100000000011101100010100010100001010000001000000000111000000001001100100100010000000001100100000000000000010101000000000011000010000001101000100000100001100011001110100100000010000100000000010000100100000000001000100000010000000010011100000001000000000001001100100001101100000110010100001001110010000100010100110000100000000010100000010000101010000000100001010000000000100001000110000101101110101000110010000010010100001100110011011010110001000010011001000010001011010110010010000000100000001010000010010001000000000101000000000110001010010000000000000001011001000000000000111100000000100100000001101001000100000000110100000000010100000000011000100100100000000000100000101000101001000001000100000000101010000000010100001010010000110000000010001000000100000000000000000000000100010000000101000000000010000000100000110000100000011100001000010000000000010001100100100000000010000001000000110001100011100100001001000001001111010000000011000001000000000000011101000000000001010011001101000011010000010000101000001010000110011000000010000110000000100000010010100000000010010100000100010000000110000000000100000010001100001000000100110010001100010001001011000000101000110000000000000000101001000011010101100000000000100000100000101001010100010010100101101000001011000010000011000001001101101010101000000001010000000000000011000010101010000001011000010010010001001000001001100001000000001010001000000001000010100001000000000001100010001110000100000011000001010111100010010101000100000000010000000110010100001100000001100000001010000011000000010000000000100110011000000000000000000100101001100010000000010100010010000100101100000011100000000100010010010000000001000000100101111000010100010010000000010000000010100100110000010010010001100000000100110010010000000010000001000100000010001000011100101100000001000100101110000000010000000000000010000111100000000000000001000011000000000000000010000100001111110001000001000000100000100001100011001001100010000000010001010010000011001000001000000001000001000000000000100100000001000000000101000010000010000000110000010001010000000000000101000110001000110000010001011010000000010100001001000000000000000110111000011100000000010000000111010010001001011001101000000000000001101001010000000010001001111000000000010001000000010000001000100000001000111011010001000001000001011000000010010100010010000001000100010010000000001000100000001000001110000111011000010001010000001100000011111000000000001000001000100100100100010100000100000001100101001000001000000000000000101101110001000001010100000100011100000101000000100001010010010000000000100100011000010000011010000000010000000100010000000001101010100011010000100000000001000000010010000000010000000000111010000100010101001000101010010010101000000010000001010000000000010000100000100101000001000010010000000100000100101000010100000001000100001110000000111000000000100110001010000000011000001010100100100000100000000001100000010111000001100010100000000101010000100000101010000101000100000000010000110001001010000011001000001000000100000000010000010100000100000001010000000100000000000010000000000000001100010111100000100001000001000001000001100000000010000100000010000000001111000011001100000000000010100001111011100100101001110010000000001001010100101100001010011000000000000100001001001000000011001000000010000010000010000000101000010001000110100000100011100100100000000010100010111001000101010000010001000000001001001000110001010111000000110000000000000001101100010000100100000000001000010010011000000000000000110000000000001010010100011100100011000000010000000001000101100000100101010001001100000001000000001011000011100010000000000101000000100000010000010000000100101000100000010010100001000000000100101001000100000011001000000010000100000000000000000000110100000000000010001110000000101100000011000010000101000000000101011111000000000010000010001000111010100010000001100110001000100011000010000010000000100000000000010000010010011100000011101000101000000000010001010001011000000000100001001000000000110000000101100000010001000000000010000010001000000101000110010001000000110001000000001101000100000001000000000101111100001010000001001100000000000001000000100000000001110010000100010001010100100000011010000000010010001000010000100000101101010111010010111011000000100010100000001010000000001001110011000000000100000000001100000100001100000000001010101001011000001000110001100010000010000000010000011100000000010100000100100010000000101000110000001100001100010000001100100100100101000000001100001000001100000100000001100000001000101001000001000100101000000100000000100000000100010000011110010100001000000010100000001010000001100100010001001000000100001000001100000101001001000001000000000101010010001000010110010000000011000001110010001000001100000110000001100010000000101000010111000001000000010000000110010101010011000000011000010000000101000100100011000000000100000001000010100100000000010000001000000101010000000000100001000011100001000000000000100001000000000000011110000001000000100000010110111100010000100000111000000000101110000001000001001110000100101001001100000110010000001000001000010000011100000000000101001010010100001010110000100100000011101100000000000000001101110100100",
	"1111000011010000001100000000100010100101000000011100011001010000000001000000001010001000000101110100011010010000001000100000000101010001000100110000010000010010000000000000100011010100001000001001000100000001001100001000000001000100000001100111111100001000010000000001101000001101010000100011010001000001001101000000010000000000000111000000001100001001000000001000001000000000010001010010000000000000011100011101000001010001011110111000001101000110011000001010000000000000101000001101000000000101100000100000000000001000010010101010000000010111011000100100101100011000000000000001000010000000000100000000010100010000000111110000100000000011000000010001000010010101110000000010000000001000110100000100001100000100010000000011001100000000101100001011010010001000001011000000110000111000011000000000001101000101101110110100101110000001010000000100000110000010000000100000000100000010100000100100101010000011010000010100001000100001000101001000011010001000100000000101110000000100000111101001011010101100000000001000000000010101000001100000010001000110100001000010101100000000000111000000110100000100010000111010001001010110010000010000000101111001001010000001100010100000010101010010000011000000101000100001010000100100110101101000100000001010010000000011000000001000010000010010110000011001011001000100110001000100000010000111010100001100000000010010010000001010000000000001010000000001000001100000001100110101100000011100000100000000001000001000000000000100011000110001000001000000000000010000000000001100110011101000001000100001100000001010010010000000110100101000000000000010100000010010000000011010100100100101100000000001000010100000011000001010110100010000100000110010000000100010100000110100101000010110000000000010110001100100000000000000100100000000000010101000000001011010011000010000011000000001000000000001001010001100000100000010000000000101100101001000001000100010000000001101001100101010100100010010001010000101101000001000101000000110000000000000010000010000000010000000100001010001000001000010010000000100000100010000000000000000000001100000011100000001100001100000010011110011010000100000000000000000000000101100000010000000100000000000000100000100100001010100001100011000010000100000101100000001001000011000001100010100010000000000000001010011010000100000110010000010000000001011010110000010100000000000010001100100000100001100010000010000010110000010110010010001100111011101000000011000010000110010000000000001100000000101000001010000001100000100100101100000000000100100000100001000000110000000000110001001000111000100000000000010100000001000001100101011100011100010100110111011000001000101000001001000010000000000100000001000000100010100000000101110001100011000111000000000000001110100010100010011001000010010000000110110000010000010011000000001000001010011000000000001011111000000100100000001000101000000000101011000000000000001000100000000101100000001000000000000001001000000001000000000111001100110000000001000100100001000100100010000001110100101100100001010101110100100000000100000101000001000100101110011000100001000000101000011010101010000001100100000001001000010000000111111000010000010011000000010000001100101100001011000001001000001100010101000100010100010000101100010001001000010000111100100000110111101000100000001111000000001001001010000010001000001000100000000000000101110000001000100100000001000100100010101010100010001010010010010011000000001010001011000010010000000000000000010000100000001010000010110010000100000000110000100000100101001001101000001011010010000101000001000100011000010100001100000101010100100100001010000001001000011100100000000000000100000000111000001010000000100000000000010010010000001000000000010100001101000010100000001000110000100000000010010001010000000010001100000000011001000101101011010000000111011000001001010000100010000000111101000000100001000001000000010010001010000000010001110010000001011000001110000000000101100000000101000001000001011000010000100000000010000101000100000000001001000100000001000000010000000000101010000010100000000010010010000000100010001100100100001110000010000000001000001000000010111101001001010101000001001001001010001000000001100010100000000010000001000110001000000010000010100000000000100000010001000101101000000110000000000001000000000000011000000110000001000000100000011000011001001010000010000100001001000011001010100000001000001010000000110000111101000100110000000100101010110000001101000000001010001010011000000010000010110000000000001000011000000010010100010000000000001001000000100110000001010000001001010000000100000000101000000000010000000000001000100110100000011000100000000000001000000000011011001010001000010100000000000010000100110000010001000000110110000000100001100010000010000100100010010101100001000010100010001000010100000011000000000011000000000010110000010001100010010001100000100000000000000000000000110000000000010000000100110000001001100011000100000100010000000010001111111100000001001100000000000000000001000100000010000000000101000100001000000000101000111000101000011000100001101110100100100000011100000010010000000010000000000001010000011000000000001100110010100011000001001100100101001000001110111000011001100000001100011110100100000000110010100000010001000000100100110011011011001010000000100110010101000110000001011001001110110110101000010000011000000100000000011001000000001010010010010101100000100000000010000100000001000011000001001000001100000000000001001000000001100001000010000000100101001011100100000001100000000010001110000000000000001100000000010100110100001000010000000000001000100000010001000100001000101001010000001100001000110100000001000110001000110110001001000000000100001100000000000011010000010000010000100000010000010000010100101000000010000010000000000010001000001010000101010000010100000000100000000000100001100111010000000010000000000110000000010111000010101011010001000000010001010010000001001000111010000010010000000011000110110010000000000000110010000000001000101100101100000101000000000100000001101100001000100100111001000001010001101001001000101010000000000000010000010000110101100101100000100000000000100100001011010000010100000100001000000011100110000000000000100101111110000001000000010000100001001011010000000010001001101101010000001010010000001010000001001000100000000010000000000011000001000001000101100000000000010111000001000010000001110000000001010111001100110000001110010100000000000000000000001000000001000000001001000001000100011101000001001001001100001000000010000000000010000010000000101000000000000000000100010011011000000011000000100000100001010100110000000010010100000010000010110000010110000001100000000000000000110010011100000011000000001000111000011110000000010001000000101010000000001011000000010000000111100010010010100000000001001000010001000010001111001010110000000001100011101000010000100111000000100010000001010000111010001010011010100000101000010001100000100000100000000100100100000000000000110010000000010000000100110001000000000100000100011100000000000001010000000000110010011000110001100001000100100000010100001000000000000010011010000001001100000000000010100000100000010010000010100001011000000100010100001000000001101000100010100100110110000101010000000001001000000000111101010111000001000101011100000000000100100001001000101100000001111000000000110100001000000011100000000010000000110000110001000100000100000101001000010110001000000000101000101010001001100010000010110101000000000100000100000000000010010000010000000100000000010100100100110010100101010010000100000000000001100010100010010000000000010100000000010011110000000000010100001000001001000100000010101010010000001000100101000100100100000000000000001001000110000000000001000001000000000000000001000101000000000101010000110000110010001110010000000000000010001000000010100101110101000000000001000000000011000000100010100000100111010001100001101001000000000000010000100110010011010000000001001100101111000000010000010000010000000000001001001000110100000000101010000010001000000000010010000100100100100001010110000001000000000010000100001010100010000100100100000000100000001000000001100000110000000000001000000100000000101000001100101001000000100000010000001011001000000010101000000000010010000110000000000010000110000110100000101000010100010110000110000110101000000110010000010011000000000000011000010000010111000000000100001010100000001100000010100000000001001000000110001000000000000000100100000001001011100110000100000000000000010100010101000001000000000101000011001000000001001000000010000011000000000000001100110011100101010000010000010100110000100100010000000000000010100100000101000001000010100010000000100100100000100010001000100100110000000100001111001000001110100011001010000100001000010111100110000100000000100000011000001011000000000000100110000000101010110011010000100000001000000101000000000001001111100001000001111010000100000000001011011000100000100010001000000000110010000100100000000011000000001001000000001000101100001010010000100000101101000010000100010000000011000000100100011100001011000001000100000001000001110010100001001011010010000000101000000001100000001100000010011001010000000101000000100100000101000010100011001000100010100000001000010010001000111101101010000100000000101000000010001100000011000010001001010000001100100001110000001010000001000000101000000010111100000000000010000010000000001011000000001100000001001010100100100100000000001100001000001010101100010101000010001010101010000000000000100000000000000000101000000000011000011000111000010000101000000000001010111000001000110101000000000100001000001100000000001001010001001000000101000111000000010000010000000001001001010100000000000000010000001000100011001010101000010001100000001000011010100011000001100001001100011001010100000001000000000011000001100101001101000000001111000000010000000100100000010001100010100001000011100000000000100100010100000000000010010000000001001110001000011011110100000000100110010001000110111101010010110001000000000100011000000110000000010000000000001100010100000110000000100101000010000100000010011000001010001110100100111000000000001000011010000",
	"0011010001000010001100000000100010001100100000001000011000110100000110000001001010000001000000100100001110011000000100100001001101010111100001111000011000010001000110000101100010001000011011001000000110000000001010001000000110000000001001100001111000001000010100000001100000001100100000101011111001001110001001001010011000001000000110100001001100000001000010110000000010110000010000011010001000000110011000000100000111110101110100010001001001010111000000001100010001001000101001001000000000100101101001101000000000000100010010100010000000100110110000100000000100001001001101000001000000001000100100000000010000000000001100101000000000010001000001010000000000010100110000110110000000001000011001100100000010101000000000001011000100000010110001000001110000100000101011000000000000011010010000000010100011001001100000000001101011010100001001010000000100101000000110000000000000010010000000000000101011110010000000000100001000101100000100111000001010010010101100100101100110100001100110001001011010000001000000000100100000000101001000111000010011111010100001100000101110011001101001010000111100010101001000101010001001010110010000000000010001010001001110000001000000000000010111000010000000000001000010000010000010100101001101000000100100001000010000100010010000100000010000000000100110110001001001001100110001110010000010001010000100000101000101000000000000001010010001001001000001110001000000000000000000010000001000011010010100100010001010001010010000000000011001001000000000010100000000110000000100001000100010100001000010100100100000001010000000001000111100001000100010000000000000000000001000010000000010100011000100010000000100100001001000001010110000010000100000100000110000001000000000110100000000010000000101001100101001101101000000000001110000000000000011000011000000000010011001000000000000001001000110100101010000000100001001000010100101000100010000001100000000100110010000010101010100011000000000110010001100000001001101000001100000000010010010000000011011010000001010000000100001000000000001000000001000000000101000001001000101011000000000010010000000010000100000100000000100001011000100100000011001000000100000101000000011000100000001010000110101100010011000001100101000001010011001100000101000100001011010011000001001000100010000100000001000001011000000100000110000000000010010001010000010100011100010000000110000110110000101001001000010010001000110000010000010010000001010011100100011111001010000010000010001001001000000001000000000100000001000000000000100010000011000111100000100010000000000000000000101000010000101100101000000101010100000000000000110010011000011100110000110111111010100000101000001000000000000000001000001000000000111000100010000001001000000000001011000000000001000000101000101010010011000001010101000001000000001001010010000100000011000100110100000110000011111000000000000011001000000100010000101000001100000100101000000001000000010010000010101000001001001000000011000000100101000100010000010100000000000000110000100000000001100000110110101001000000110100011000000110001101100111000000101100011000100001000000101000010001000100100000100100000010001000010000000001111000010011010011000000110000001000001101101011000001001001001000110100000000110101011000100100000100001000001101100100110011011011101001100000001011000000000001000010000100000000101000000010001000001101001000001000000000000100010110100010101100101110001111000010100010001000000100000011000001000010000010110000010000100000101000100110010010000000000000110000110000100001001000000000000000000000101100000111010000001000110000000110000110000110000100000011100000000000100100100010000000000000000000010100001010100101000000100000000000000000001011000000111100011000011010110010001000011100000010000001000100000000100100000010010010001000000000001001010000000101010100000100100001000000000001100100000100000000010001100000000011000001000100010000110010100000011000001010000000000101000001000111000000000001011000000010000001010000010111000101000000010000000000000001010000010000000011000010000010000000000010100010100100001000001000010100000010000011000000011000100000010100000000001100010101000010100001000101001000000000000010000000000000010001000000000000100000000011000000000000100000000101000010001000100100000000000001001000000010011000101010010011010000000000011001011001001010011010000100001000000000000011110000011000000010000000100000011101000000110001001100101011000010000101000001001010001010001000000000000110010000100001001000010000000000010110010101010010000000000000011010100011010010001000000000000001000100101110100000010000010000000000100110000000000000000001000000000000101000011001101010001000110000000000100010000110110000000000001000110000010100001001000111000111000100001010001000010011001111000100011000000100100011010000000011001000001010011000011000010000000000100100100010000110000000100100101001000000010000000100101010010100101011100000100101000000101010001111000000000101001100100100100100000001100100000000000000010000000100111010000000001001011000000100101101100001101110000111000010011000000001001000100100000000010001110000001001010000001000010001100011001001001100011101101100000110111000000000010000001101010100110001000010010001001000010000100010000100000001011000000000100001010110000001101000100010110011000001010001000100110001010010100000000010001001010000001011110010000111000010100000000010000010000001000010000001010000001010000000110001011100010100010001000010100110100100011011100000000000101001010000000010010000000100010100000000010110010100000100000010000000100000000000010001100100000100001001010000011000001000101001110000011110100001010010000010000000001100001100110000000000000000000010010100101000100000000000010110110000010010010010000000100000001000001100100100010000100001001011100100001000100001101001010000010011000100000100000001001010000000101001010011000001010010000011110000000010111010000010101000000100010110100010000000000000110000000010010000001110111000000100000000000100000000101100000000000000000011101101010000000011000000100000010000000000000000010001110001111101000010000001101000100000100001010000010110000100001100000011101000000000010001001100011001100001000100110000100001000011010010000000001001100100010100001000001000000000101001001000100010000010011000000101000000010001000101000010000110010011000000000010010100110000000111010101001100010000001000000110011000000001101000000000000011000000000010000001100000001000000001000001001100101001000010001000000000110000000100100010000010100000000100010010001000000000000000100100100001000100110010000000110100000000100100110000001010010000110000000100100000100010011010000010000100000110010000011110110000010011000100101010000000001001000000000010000101010010000100000011001010001000000000000001000010001110110001000000100000001000000000000101011000100000000011000001011010001000111010000000100000000001000000100000000100011100101100000010001000010010000000000111010001001001000000000101000010000000000000010000001000000000100100111000000001000000000010010000000100000000010001000111110000001001001101000100000011000000000101000010000010101001010000000000000100001000000001001000000010001110000000001000010001000000001000100010101101010111000101000101011000011000001100100001011000100000000010111100000000010100000010000011101010001000000000010100110000001110010100000001011000010000001000000000100000100001011000100010000011110001000000011100000000000100010001000000010000000100001000001110110110001000100000010000000100011000000001100010100010010000100000010000000000010001000001100000011011001010011000010000001000100000000000101100100111000000110100000000000000100000100010010001000001011001000100000000011000000001000000000100101010000001111000000010100011001100000000010000000100110001101001100000100001100000010000000100000000100000000101010000010000001011000101100000001000000100100100100010000010001000001011000000000000000000000000000100000000011001000100000101001010000110000000001100000110000100000101100000010010000000000000000010100100000010110000001001000000011100000000000000100000100010110000001001000000100100011000011100111100101101001001001000010100101000000000000000000000000010010000010100000000001010010110010100001001000010110001000010110110010000001000100110010000110001010000000001001000101000010101000100110101001000110000100100000010100110000001001000000010001001001101010000010100000101101000000011001101000010000000110000010101000100000000010000000110001010000000000000000010100010000110000001000100011011000000010100000000000010010000100100010010100001010000000000100011010101000000100010000000100100001010000000001000110000110000000100000010001000100110100001100000000101000000000001101011000100000000000000011100110011000010000011000010000000101001000001000000000001000000000101110001011010000001000011101001111011100100010000010001000000001000000010011000000000001101000101110000000011000000000011000000000000001001100110000001100000101101100010001101000001000101110000000100011100000000100000010000000001000001111100100001000000110000000000011000000001000000101000000010001000000000000101100000000001010110010000000011000110000010000100001010010010000001011100100011000000000000111100000011000010011000011010010101011000001101000000100110001010000001000000011100010010111100100000100000000010000000110010010100010000000001000010100000101101000000001001000000001100000000000101010000001010000000000000000100100000000000000000000000000100010001011000010000011000110010100000000000010000101100001101001000000000000000001010000000001001000000001000000001000010000000000110010000000010101001110110001000100100001110001001000111001010111100000101000100001010001010100010010100100010000000001001010010000000000100100010000101000010001100000010100000000000010000001000000101010001000010001000100010100001001010100101110101000000000010011100000000100010000100001010001100010001010100100100010110010100010010010000001100000100000000001000000111010000011001001000010101010100000000100000001010010000101000100000000010001011101000101000100000001001101100000",
	"1101010000010010001100000100100011111111110001011000011000000100100010000000001000000100010101110100100010011001001100000010000010100111011000011010001010010010000010000101000001011000001010000011010000000001001000001000100001010100101000000111001100101000000000000001000000000000001000100001111000110110101001000110010000000000001111100011000100001000000010100000001100010000110000001010001000000000000100001001000011000000001000001000101010010111010001001100010001001000011001100001000100100100101001000000000000001000001010100101000000111110111000000100101000010000001001000001000110001000110100000100000000000000000100011000100000010000001100000000000010000000100000000000000000001001111111000100001110101000010000000001000000000000010000001011110010101000110010000100010001110010001000000001000010010001001110101100000001001101000101011101001110100011000011100010000100000000010001100100101001100010000000000101001100100000000000001000000000101010101000000100110000101000000001100011011010001101100001000101100000100000001000100001011111111100100010000010100101001000101101010000100100011101010000010010001100000010010100010000001101011000010000000000101000100000000100000001000000000101101100100101110110000101101111101010010100000000010000100010011000101000000000010001000110111000110001000100010000010010000010011110010000101001000000010000000000000010010001000001000000010001000000100000000100000000100000001110100100100000000010001000010000000000011100011001000001000000000000110100100000001000100000001000010010100000000000000010100110000000111100101000101010000000001000110000000010001000100000100001010110010001000110100001011100011010100000011001000000000001110000000010100000010100100000100000100000000000011000000000000000000011000100000000000011101001000000001000001001001000001000000000010100000011011010000101001001000010100101000001100101001100000011000111001000010101100100010010101000010010010011000110001101000010101000000100100000000000011011011000000000000000001000000001000000000010011000100000100001111001100000011010010001100000000000100001100000100100010010110001000000100100000101000000000000001000000001000100110000001000000100100110101011000010001100010010011010100000001100100001110010010000010000010100000100100000111101011000010010000000010010100111000000000010000110100000100100001000010000111100000001001001010010000001000000001000010010010001101111001100100001011001010000000011100001001000000000001101000001010000000100000100100000101000100000010000101000011000001110000000100010001010100110100000000000100010000000001000100000111001100011000000100110001010000101000011010001000100000000001001110101001001000110000110000000001000001000011001000000010010000001010100010100010100000000110001000000111110000100001100101000001011000000010110000000100001010111000000100010010001000101100010000101010001100000100100000110001000100100011000010001000101000001000000011010100101110000000100010000000010000100001010100100010010101100000110100101000000100100000000000000010000101100000010100001100011000000000000000000000111000000001000011100100000000000010000000000001100100010010010010000000000000101100101000001010000001000011000000110000100000110110000000001100000100000000001000111110000000000100100101100000000111000000000001001010000010100000100001100000101000101100101000001000100000000000000010000000000100000110001110010010100011001000001100001001000011010000000010010000000010000000011010000000110000010000100000010000000000100101011000101000101011001010100001000111010000010010000110001010000010010001100100000000100001000001000100100011011000000100000000010000001010000101000000000000011110110000011011011000111100011000011000110010101010110100000010000010010101100000100000001110010000110010000100101010000001000101010100000100100001101010000000010000000000110101000001000000000011001011110100011000110000100000111000001011100000100000000001000110100000010001001000000000100001010010000001100000000000010100000100000000000000010000000010000010010011000000100010110010100000000000000100110100000010000001000000011000100000010000011000001001000000000011101000000101000001000000100010100010010010000000000100001101100110000010000000000000000011010001000111001010110000001000000101001100000010011000011100000000000000100000011101000101001010011010000000000011100001100010111000001000001000000000000000101000000100000000101100100000100010000101100000001010011010000000111000001110110000101001000001000000000011001110000001110000000000000001001100000000010000001010000000000111000000100010000000000010000000100000000000110000001000100000100010100000001000010010001000000000010010000100100010000010010000001000010000100110010100001001111101000111000100101000011100110001000010100000011000000000100000000100000000001000001000011001001111100010011001000000000000000010000010100100000101001000000010000010100010001101100000100000000001010000100010001001101000010100001010000000110100000000100100000010000000000101000000100000000000101000001000100100011001100000101000110100100110000100000010000001100010000000000000100000010000000010001000010001000011001001001000011110001100000000011100010001110000001101000100110100100010110110100010000001000010100100010010011000000000000001001000000100011000001000111011000100010010000100010010000010000100000000001000000000000010000010001101000000100000011010000000010001000010000101011000000010100011011001010000000000001000000000100010110101000001000000010001001001010000000100110000000000010100010010011000100000101100110000100000101000001001000000000010000000100000100000011100001000000100100001011100001001011100000010000000101100010000110000000010000000010010000000100000010000110000011100101000100010010110010000010110000000011000000101001100000000100101010010000000000011100001000100010000000000001111010000000110000000000011000001001101010001010001000001001011100000000110001000000111000010110000000000010010110000000011010000000010101100000011000000000100100110000001001000100000101011101000010000101111000010000000110001000100000000010001110010011101100010100001100000000000100000110100010110000001100100000011011000000011110000100101111110101001000100100000000001001001010010100010001001000000011000101001011000001001000001000000100000001110010001000001100000000001100001100010001000010111000011000011010101010010010000010110000100000000001010010000001100000001100000001011000010000000011011000000000000000000000001000001001100000001100010001000010110000000000100000000000000100000000100001000010000000011001001100101000000010100010000001010010000000010110100110000010010000001110000000000100010000011110000000000001100001100011000011100111000000010000100101010000000000010010000000010000111010000001110000110100001000010000101000001000111101000000000000000100011001000010101100111011000101110000010010000110010001000001000100100001100000000000000000000100100001100010000000010000010110011000000010110000100111000000000000100000010001100010000010001011010000000110110000001000000000101000000010000001100001100000000010001000010000000001000101100000000000001100100100000000000101000100000000100010111000000000000100110000010101010111111011101010100000001000000000000000100010101010001000001010010010000001000100000010000000100000011101100000000110100000010000010000000001000001000011000000101101110010000000101010001010010000000001000000000101000100100000001000010010000100000000100010000000100010010000110000000000000101000101010110000111000000000010010000000100000000001001000000001010000100100010001100000000011000001000000010100111010011101000100001010001000000000001100000111100100110000000010010000001000100000000000000000011000000000000000111001010000100000000101010100110001011000000110000001000100000010010000001001010001000000000000010000001001010111000001000100000000000001000000010001000000000000000000000000010110110101011000000111001000000111000100001000010000000000000000001000011011000100000100101010000110011100001100010010100000000101000001000010000100000000000010100100000000000010001011010101001100100000000000100000010010110100101000000000100000000001010100011100101100010001011000000100100111000000100011001000000010010000010100000000101010000100010111101000000000010000100000010010110000100001100010010000000000010000001000011010001001000100000000110001001010111001000000010000000110100001001000010010011001000000010000010000000100001010010100110001000001000100100100000000000101100000000001010100000110000101000000000011100011000000000000001001000010100000010000010000010100011000000100000000000010010010000100101101000001000001001010000010100000000011100011000000100100110010000000001101001000000010000011000000100000000000000001110110010000000000110000001000000000000010000001100000000000000001110000110000100001101000000101010000001001001001100000001000011001100100010101010000011000001010000000010000000000010100000101110000000000100000000011000000000000001001100100000000110000111010001100000001010001000100100100100101110100100011000000011000010001000001101110100010000001000000000100000000000000100001010000000000000000010000000001000001100101000101000000101011000100100000100000000000010010000000100000000010000100000000001110000000001010011010001010001100010000000001000001011110001000000000000000110000000010110100100000110010000000001000100011010000011100100000000110100100110000000000000001011000001110101000000001000010001010100000100001000010100000000100000000000000000000000001001110100000001000010000000010001010001001000000100101001000000001000000000000000101000001000000011000000100011001000001011010000000000001100001111010001000100000000010000000000111001000110001000001100100100010010000100010000100000010000100011001010000010100000100000000001010000010000001100010100011000000000000000000100000010000100010001001100010000000000010000001010001000000000000010000000001111100001000011111000000010000100110110000000110101000010010100000001100000000111101000100100000000000011001001100101100010010000000000101001010000000000010101000001000001100101100110000100000001000000110010"
	); 
  	variable actual : testactual := (0,1,2,3,4,5); -- this is an array of what should really be predicted (first test should be predicted as 1, second as 0, etc.)
	variable numtests : integer := 6; --number of test inputs we are using
	variable correct : integer := 0; --counts number of correct predictions
	variable total : integer:= 0; -- counts total number of predictions (i guess this is pointless, we already have number of tests we are running)
  begin
	for i in 0 to numtests-1 loop
    		result <= classification(test(i), testclasses);  -- calls function given a test input and the class HVs
		wait for 10 ns;
		if (result = actual(i)) then --checks if result from that function call is equal to the actual class of the test input
			correct := correct + 1;
			total := total + 1;
		else
			total := total + 1;
		end if;
	end loop;

    	wait for 10 ns;
    wait;
  end process;  
   
end behave;