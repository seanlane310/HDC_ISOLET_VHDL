library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity declarations is
	PORT( A : in  STD_LOGIC_VECTOR(31 downto 0);
		counta : out STD_LOGIC_VECTOR(15 downto 0));
end declarations;

architecture Counter of declarations is

begin 

process(A)
variable count : unsigned(15 downto 0) := "0000000000000000";
variable B : unsigned(999 downto 0) := "1011001101001111101111011001000100001110100000101000110011000111111010111011111101011010100100001110000111110001000001000010011011100110010011001011100110110001110000100011110101101100101010001011111100000100111001101100010110101110001111001101110101010000011101110001011111000100101110010011011101101110101110110110010010001100010010001100111100110101110011101111111100111101101010000011111000011110001100001011100010101001101100011010111110000110100011100111010101101000001000001111010111111110011101001010110100111101111111001001111000110101110011111001000010110100111001000010001110110100011100110110100000110010001010110111101111101001000100000111111110100001101010100110101010101101010101101010001111011001101011001000010110001111010000111001011100101110011010110100000101101011101110011010110000000101001100110100101010011110111100100001000111111110010110001111011100100011101111010010011011101100101010101101001001001101111000011010111101001100101011101001110111010111101101010001001100100011";
begin
	count := "0000000000000000";
	for i in 0 to 999 loop
		if(B(i) = '1') then
			count := count + "1";
		end if;
	end loop;
	counta <= std_logic_vector(count);
end process;

end Counter;
