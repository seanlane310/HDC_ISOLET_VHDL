library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
 
entity testing is
end testing;
 
architecture behave of testing is
 

	type slv_arrayclass is array (0 to 5) of std_logic_vector(9999 downto 0); -- length of this array must be number of classes (letters) we are tested, vector length is dimensions used
	type testarray is array (0 to 5) of std_logic_vector(9999 downto 0); --length of this array must be number of test inputs we are running
	type testactual is array (0 to 5) of integer; --length of this array must be number of test inputs we are running
	type samearray is array (0 to 5) of integer; --length of this array must be number of classes we are using
  	signal result : integer;
  	--signal total : integer;
  	--signal correct : integer;

  function classification(
    testinput : in std_logic_vector(9999 downto 0);
    classes : in slv_arrayclass)
    return integer is
    variable closest: integer:= 0;
    variable mostsame: integer:= 0;
    variable numclasses: integer:= 6; --number of classes (letters) we are checking
    variable numdimensions: integer:= 10000; --number of dimensions for HVs
    variable same: std_logic;
    variable amountsame : samearray := (0, 0, 0, 0, 0, 0); 
  begin

  	L1: for i in 0 to numclasses-1 loop
		L2: for j in 0 to numdimensions-1 loop
  			same := testinput(j) xnor classes(i)(j);
			if (same = '1') then
				amountsame(i) := amountsame(i) + 1;
			end if;
		end loop L2;
		if (amountsame(i) > mostsame) then
			mostsame := amountsame(i);
			closest := i;	
		end if;
  	end loop L1;
    return closest;
  end; 
   
begin
 
  process is
-- store classes in test class array 
-- store test inputs in test as an array of test inputs
-- store the actual value of the test (whether a,b,c,etc.) in testactual array
-- store number of tests you are conducting in numtests
-- loop will run tests with each of test inputs to find what class it most closely matches
-- it will return that index as result
-- if index matches the actual expected result index, correct counter is incremented
-- the total number of tests conducted is incremented regardless of correct or incorrect prediction
 	variable testclasses : slv_arrayclass := ("0000001101001101101110100110000100101001100000100000000000001011111100011001000000000100110001000010110111000000010001101011011000000000100000000010110000010101000000100110110000011111000000010000000000000111111000000100000000011000000000000011000010000000000001011100000001000001011010110000001111100001010110010001110000000000010000001110101100000010000100000001010101000000101001000000001100000001101000100011111000001011011001110010010101000000000100000000110001110000000000000000010100110001000000001010110110110000100000100001100000001111100000001000000000100000100010010000010010000000000000000000000000000000000100111000010000000101000000001010010001010010010100000000100001100000000001100000001000000000100001000000010100111100001010000000000000000101100000000011010000000011011000011100001001101100000000000000000010101010101001001100011010000001010011000001000000010000000100010000001000000000001000000000010011011100000011100010010000001110010000000000100000011000000000100000000101100010001001101000010000010100100000100000100000000011110000000000000001000111110000110100100000000000000000011100000000001011010000011110000000000101101000000001000000000011111010000010100101110000110000000000101000000100101100000111000111000000010000000001000000001100100000000100000000101100001110101111100011100000000000100000000000001000000000001110000100001111000100000110000000000000010000000110000000000000000100000100000000000101011000000000000000010000000000100101000000110100000000001100101000000000111000101011000001101000000000111100100010000010100001000000000100011100000110110001111100000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000001000001010010000100110100000000000000000000011001100001100000000000000000000011000000000001100000000000010000000000110010000000000000100010000000000111000000000110000010000000011100000000000100000010000011000000001010110000011000110000000000001101010000010000000100110000000000100000001001000000000000110001011111011100000000001000010011000000000000010111000000100101000000000000000001100000000100000001000000000000110100001000101100111101100111100001011001100000000111101001110111001101000100010000000000000001100000011000100000000110000010000000100000010100000000110000000000100010000010100100100000000100000000000010100000001000000100010000000011000000000110000011001000101010100000010101001010000000000000000011100110001011110000001111001010101101000101000011111100001100010110000000000001101000000000000000001101000100000000000000000011100110110000000000001000000001011000100011100000110000000101000001011000000000000000011010010001011000010100101100000110000000000001000001000100000010000000000010100000100000011110001000000000000100011100011111000110000110010000001010000000000000000000011000100100100000011100110000000001100101001111010111000000000000000100000000101100001011111000000000011000010010100000000000000111100001011101100101100000010000000000111110000000000000001000001000000000000000000101000001010000000100001000000000011000000111000110100110111000000100011010100001000010110010000000101100000101000001000000000100000010000001011100000111001100000001110011000100000110000111100000011100001000001101010100000110000011111000000010110000000001010101010100000101000010001000100000001100000000001000000100000000000000010000001101100011001100001000000000000100000010011111100001100110001100000100001011101010111000000000000001100000100100000000000000001100001100000000000111100011000000101111010110000000010011000100000010000000000010000100000001000011000000000000000000000001001111010000000000000011101100000000001100000000010000001000000000100000000000000001110000000000000000010111000000001010000000111010001110110000000000111100100000000000010110000001000000000100010000000000000101100000000001011001101110010100000000000100000000000001011010001111111001101001011000001111001110000100001001110001001001101001000011100000000000000101001000010000110010000110101001000000001000101010000000000000000000111000111010100100100000000000010000000000001010111000010000101011100100000000010011000000000100101000001101110000000000011100000000000000000000000000101000001111000001100000001101101001001000100100001011010111101001000000110000100000000000011100101000000000000000000000000000000000000000000010001001100001001111100011000000111000000000010011000000000000000000000010000000000010000000000001110110000000000010000000010100000000000000000001111101100100000000000001000000010000001000000110010000000000000000000000110000000001000110001010010010000000001100000010101011110010100010100000001001001100000000000000001101101000001100000011010111011100111000010000001101011011000000010000000000000000000011000100000000000000000001000001110000100110110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000011000000000000010001100001110011000000000000000010100000000001000111111000000000000000000010000010100110110100000010100010011110000000110000100001000000000000100000000100000001110010001011100000000000100000000101000000010100010101010000000100110100011000100000000001001011100001111100001001010000000000001000000000000001010000000000010010110000000111001111101001101101011011000000000000111100000000110000000001011000000000001000000001100100000000011100001100000010011000000000001110010000010010000000011000000010100000000000010001011100000001101100011110111010011100000000100110100101000000010001010000000001110000101101101001100011100000000110001000000000010000000010010011010000000001110000000000000000001000000011011100000101100000000100100100010010000000000110000000101110000000110000011111101110000000001011100000101001000100000000010100000101000000100110101000000000000000000010000000000100000001111000001101000001100000001000010000100000110000000010111010001011001001000000000100000100100100000110000101011000000000011111000000000000000000000010110100000001000110000000000000000000001110000100000000000001000000111010000110000101101100101110000001101011000000011111000111101100100010000001000000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000011110000000111100100000000000001010010000000110000001000001100001000011000000010000100001000000000001100011000000100000101010000000011010000100000111000110001000000001001010110010000100110100010000000000001000000000100001000110000101110101110100000000000101000000101000001100000000001100010100100100000110000000000000000010000111001000010010011000000001100000001100000100000010010001101001010010000001000000000010111000000100000010000000000001010000100110001100001100011000000001111000011000011000000001101000001010100000000000000110010100010001100000001100000000001010010000000000000000001000001110011111000010100001000000111100000000001000001010000100000000011100101001111010000001001000000000111010001100001001010001100000000000000000000000000001100010000000000000000011000110001100100100001000011000000000001001000011000001000000000110000000000000000000000000011011000000000000000000001000000111100000010010100000010011100000001000001101111111000011100010000000000000100000000100100000001000000000001010000000011000000000110111100000010000000000100101000111010001000000000100000000011010100000011100000000010000000001010000000100000110000100000000011000010000000001000000010000010000011010000000000100000110000110101011100100001110000100100000010101000000100000000010000000000000000000000000000000000100000001100000110011100000000000010010000000100000110000001000110000001100110000000000100000000100110001000000000001110010000000000001000010010111001100000000101111011000000011101000001011000000111100000000000110000110010000100001111011001001100000011000000000011100000000000000000110000010010000100000000000000000110010010001000001000000000011001000011100000100000010100000101100000000000000000101010000011000000000011000000000111001100000000000000010010111111110000000001011000000000000000000001000010000000000000000000000010000101000000010110010000000000000010101101110000001101000000111010000011100000000001100000000100001011000000110000000000000000000000000000010000000101000000000110000110010000000000000000111001000111000010000001110000000000000000100001010000000000000001011001100000000101111011100000000000100001110100000100110000010110000010111110010100000000101100001001100000000000000000000001000110000110001011010010000010010100000000000101001110000000000000000000000000000001010110001100110100011100100100000000100000000000101000011011010110000000000100011100001110100000010000110011111110000000010110000000000000000010000000000000000101010000100001000010011000100100000010010110110001111110101000000000000000000010100000100011010000001000000000000000101000110000010000100100100000001010101111000000000000000100000101100000001011000000000000000001010001001001010100000001000000000000001001110101110101000010100001001010010000000000010000000001001000000000000000000110100000111000000010101111100000100101111110101110100000000111010000001000000001010110000001100000000000010001010010000000001110100000000001000000000001101010100001010000010000101010100110101000001010111010000000001100110000000000000010000010100000000000010000000000010000000000000000000000000000000101100000001000100011100010001000011000000000000000000000011110000000111110000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000100110001101001100000111000000011000000000000000011100000000001000000001001001000000111101100001100000000100111011000000000000000111110110000000000100000000001100000010100011100000100000000000000000000011111100110100010000000000100011000000011100000000001010101111101100011010100000000100100011000000011010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000000100100010000001000000001000000000000000110010000000000111100000000000001100011100000010100011110010011010000000000000000000101001000000010110000010000100000000000100000000000000000010001000000000011", 
	"0000001101000101101110100110000100101001110000100000010000001011111100011001000000000100110001000010110111000000010001101011011000000000100000000010110000010101000000100110110000011111000000010000000000000111111000000100000000011000000000000011000010000000000001011100000001000001011010110000001111100001010110010000110000000000010000001110101100000010000100000001010101000000101001000000001100000001101000100011111000001011011001110010010101000000000100000000110001110000000000000000010100110001000000001010110110110000100000000001100000001111100000001000010000100000100010010000010010000000000000000000000000000000000100111000010000000101000000000010010010010010010100000000100001100000000001100000001000000000100001000000010100111100001010000000000000000101100000000011010000000011011000011100001001101100000000000000000010101010101001001100011010000001010011000001000000010000000100010000001000000000001100000000010011010100000111100010010000001110010000000000100000010000000000100000000101100010001001101000010000010100100000100000100000000011110000000000000001000111110000110100100000000000000000011100000000001011010000011110000000000101101000000001000000000011111010000010100101110000110000000000101000000100001100000111000111000000010000000000000000001100100000000100000000101100001110101111100011100000000000100000000000001000000000001110000000001110000000000100000000000000010000000110000000000000000100000000000000000101011000000000000000010000000000100101000000110100000000001100101000000000111000101011000001101000000000111100100010000010000001000000000100011100000110110001111100000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000000000001010010000100110100000000000000000000011001100001100000000000000000000011000000000001100000000000010000000000110010000000000000100010000000000111000000000110000010000000011100000000000100000010000011010000001010110000011000110000000000001101010000010000000100110000000000100000001001000000000000100001011111011100000000000000010011000000000000010111000000100101000000000000000001100000000100000000000000000100110000001000101100111101100111100001011001100000000101101001110011001101000100010000000000000001100000011000100000100110000010000000100000010100000000100000000000100010000010100100100000000100000000000010100000001000000100010000000011000000000110000011001100101010100000010101001010000000000000000011100110001011110000001111001010101101000101000011111100000100010110000000000001101000000000000000001101000100000000000000000011100110110000000000001000000001011000100011100000110000000101000001011000000000000000011010010001011000010100101100000110000000000001000001000100000010000000000010100000100000011110001000000000000100011100011111000110000110010000001010000000000000000000011000100100100000011100110000000001100101001111010111000000000000000100000000101100001011111000000000011001010010100000000000000111100001011101100101100000010000000000111110000000000000001000001000000000000000000101000001010000000100001000000000011000000111000110110110111000000100011010100001000010110010000000001100000101000001000000000000000010000000011100000111001100000001110011000100000110000111100000011100001000001101010100000110000011111000000010110000000001010101010100000101000010001000100000001100000000001000000100000000000000010000001101100011001100001000000000000100000000011111100001100110001100000110001011101010111000000000000001100000100110000000000000001100001100000000000111100011000000101111010110000000010011000100000010000000000010000100000001000011000000000000000000000001001111010000000000000011101100100000001100000000010000001000000000100000000000000001110000000000000000010111000000001010000000111010001110110000000000011100100000000000010110000001000000000100010000000000000101100000000001011001101110010100000000000100000100000001011010001111111001101001011000001111001110000100001001100001001001101001000011100000000000000101001000010000110010000110101001000000001000101010000000000000000000111000111010100100100000000000010000000000001010111000010000101011100100000000000011000000000100101000001101110000000000011100000000010000000000000000101000001111000001100000001101101001001000100100001011010111101001000000110000100000000000011100101000000000000000100000000000000000000000000010001000100001001111100011000000011000000000010011000000000000000000000010000000000000000000000001110110000000000010000000010100000000000000000001111101100100000000000001000000010000001000000110010000000000000000000000110000000001000110001010010010000000001100000010101011110010100010100000001001001100000000000000001101101000001100000011010111011100111000010000001101011011100000010000000000000000000011000100000000000000000001000001110000100110110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000011000000000000010001100001110011000000000000000010100000000001000111111000000000000000000010000010100110110100000010100010011110000000110000100001000000000000100000000100000001110010001011100000000000100000000101000100010100010101010000000100110100011000100000000001001011100001111100001000010000000000001000000000000001010000000000010010110000000111001111101001101101011011000000000000111100000000110000000001011000000000001000100001100100000000011100001100000010011000000000001100010000010010000010011000000000100000000000010001011100000001101100011110111010011100000000100110100101000000100001010000000001110000101101101001100011100000000100001000000000010000000010010011010000000000110000000000000000001000000011011100000101100000000100100100010010000000000110010000101110000000110000011111101110000000001011100000101001000100000000010100000001000000100110101000000000000000000010000000000100000001111000001101000001100000001000010000000000110000000010111010001011011000000000000000000100100100000110000101011000000000011111000000000000000000000010110100000001000110000000000000000000001100000100000000000001000000111010000110000111101100101110000001101011000000011111000111101100100010000001000000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000011110000000111100100100000000001010010000000110000000000001100001000011000000010000100001000000000001100011000010100000101010000000011010000100000111000110011000000001001010110010000101110100010000000000001000000000100001000110000101110101110100000000000101000000101000001100000000001100010100100100000100000000000000000010000011001000010010011000000001100000001100000100000010010001101001010010000001000000000010111000000000000010000000000001010000000110001100001100011000000001111000011000011000000001101000001000100000000000000110010100010001100000001100000000001010010000000000000000001000001100011111000010100001000000111100000000001000001010000100000000011100101001111010000001001000000000111010001100001001010101100000000000000000000000000001100010000000000000000011000110001100000000101000011000000000001001000011000001000000100110000000000000000000000000011011000000000000000000001000000111100000010010100000010011100000001000001101111111000011100010000000000000100000000100100000001000000000001010000000010000000000110111100100010000000000100101001111010001000000000100000000011010100000011100000000010000000001010000000100000110000100000000011000010000001001000001010000010001011010000000000100000110000110101011100100001110000100100100010101000000100000000010000000000000000000000000000000000100000001100000110011100000000000010010000000100000110000001000110000001100110000000000100000000100110001000000000001110010000000000001000010010111001100000000101111011000000011101000001011000000111100000000000111000110010000100001111011101001100000011000000000011100000000000000001110000010010000100000000000000000110010010001000001000000000011001000011100000100000010100000101100000000000000000101010000011000000000011000000000111001100000000000000010010111111110000000001011000000000000000000001000010000000000000000000000010000101000000010110010000000000000010101111110000001101000000111010000011100000000001100000000100001011000000110000000000000000000000000000010000000101000000000110000110010000000000000000111001000111000010000001110000000000000000100001010000000000000001011001100000000101111011100000000000100001110100000100110000010110000010111110010100000001101100001001100000000000000000000001010110000110001011010010000010010000000000000101001110000000000000000000000000000001010110001100110100011100100100000000100000000000101000001011010110000000000100011100001110100000010000110111111110000000010110000000000000000010000000000000000101010000100001000010001000100100000010010110110001111110100000000000000010000010110000100011010000001000000000000000001000110000010000100100100000001010101111000000000000000100000101100000001011000000000000000001010001001000010100000001000000000000001001110101110101000010100001001010010000000000010000000001001000000000000000000110100000111000000010101111000000100101111110101110100000000111010000000000000001010110000001100000000000010101010010000000011110100000000001000000000001101000100001010000010000101010100110101000001010111010000000001100110000000010000010000010100000000000010000000000010000000000000000000000000000000101100000001000100011100010001000011000100000000000010000111110000000111110000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000100100001101001100000111000000011000000000000000011100000000001000000001001001000000111101100001100000000100111011000000000000000111110110000000000100000000001100000010100011100000100000000000000000000011111100110100001000000000100011010000011100000000001000101111101100011010100000000100100011000000010010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000010100100010000001000000001000000000000000110010000000000111100000000000001100011100000010100111110010011010000000000000000000101001000000010110000010000100000000000000000000000000000010001000000000011",
	"0000001101000101101110000110000100101001010000100000010000001011111100001001000000000000110001000010110111000000001001101011011000000000100000000010110000010101000000100110110000111111000000010000000000000111111000000100000000011000000000000011000010000000000101011100000001001001011010110000001111100001010111010001110000000000010010001110101100000010000100000001010101000000111001000000001100000001101000100011111000001011011001110010010101000000000000000000110101110000000000010000010010110001000000001010110110110000100000000001100000011111100000001000010000100000100010010000010010000000000000000000000000000000000100111000010000000101000000000010010010010010010100000000100001100000000001100000010000000000100000000100010100111100001010000000000000000101100000000011011000000011011000011100001001001100000000000000000010101010101001001000011000000001000011000001000000010000000100010010001000000000001100000000010011010100000111100010010000001110010000000000100000010000000000100000000101100010001010101000010000010100100000100000100000000011110000000000000001000111110000110100100000000000000000011100000000001011010000011010000000000100100000000001000000000011111010001010100101110000011000000000101000000100001100000111000111000000010000000000000000001100100000000000100000101100001110101111100011100000000000100000000000000000000000001110000000001110001000000100000000000000010000000110000000000000000100000000000000000101011000000000000001010000000000100101000000110100000000001100101000000000111000101011000001101000000000111101100010000010000001000000000100011000000110110001111100000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000000000001010010000100110100000000000000000000011001100001100000000000000000000011000000000001000000000000010000000000110010000000000000000010000000000111000000000110000010000000011100001000000100000010000001010000001010110000011000110000000001001101010000000000000100110000000000100000001001000000000000100001011111011100000000000000010011000000000000010111000000100101000000000000000001100000000100000000100000000100110000001000101100111101100111100001011001100000000101101001110011001101000100010000000000000001100000011000100000100110000010000000100000000100000000100000000000100010000010100100100000000100000000000010100000001000000100010000000011000000000010000011001000101010100000010101101010000001000000000011100010001011110000001111001010101101000101000011111100000100010110100000000001101000000000000000001101000100000000000000000011100110110000000000001000000001010000100011100000010000000101000001011000000000000000011010011001011000110100101100000110000000000001000001000100100010000000000010100100100000011110001000000000000100011000111111000110000110010000001010000000000000000000011000100100100000011100110000000001100101001111010111000000000000000100000000101100001011111000000001011001010010100000000000000111100001011101100101101000010000000000111110000000000000001000001000100000000000000101000001010000000100001000000000010000000101000100010110111000000100011010010001000010110010000000001100000101000001000000100000000010000000011100000111001100000001110011000100000110000111100000011100001000001101010100000110000011111000000010100000000001010101010100000101000010001000100000001100000000001000000100000000000000010000001101100011001100001000000000000100000000011111100001010100001100000110001011101010111000000000000011100001100110100000000000001100001100000000000111100011000000101111010110000000000011000100000010000000000010000100000000000011000100000010000000000001001111010000000000001011101100100000001100000000010000001001000000100000000000000001110000000010000000010111000000001010000000111010001110110000000000011100100000000000010110000001000000000100010000000000000101100000000001011001101110010100000000000100000100000001011010001111111001101001011000001110001110000100001001100001001001101000000011100000000000000101001100010000110000000110001001100000001000101010000000000000000000111000111011100100100010000000010000000000001010111000010000101011100100000000000011000000000100101000001101110000000000011100000000010000010000000000101000001011000101100000001101101001001000100000001001010111101001000000110000100000000000001100101000000000000000100000000000000000000000000010001010000001001111100011000000011000000000010011000000010000000000000010000000000000000000000001110110000000100010000000010100000000000000000001111101100100000000000001000000010000001000000110010000000000000000000000100000000000000110001010010010000000001100000000101011110010101010100000000000001100000000000000001101101000001100000011010111011100111000010000001101011011000000010000000000000000000011000100000000100000000001000001100000100010110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000011000000000000010001110001110010000000010000000010100000000001000111111000000000000000000010000010100110110100000010100010011110000000110000010001000100000000100000000100000001110010001011100000000000100000000101000100010100010101010000000100110100010000000000000001001011100001111000101000010000000000001000000000000001010000000000010010110000000111001111101001101101011011000000000000111100000000010000000001011000000000001000100001100100000000011100001100000000011000000000001100010000010010000010011000100000100000000000110001011100000001101100011110111010011100000000100110100101000000100000010000000001110000101101101001100111100000000110001000000000010000000010010011010000000000110000000000000000001000000011011101000101100000000100100100010010000000000110010000111110000000100101011111101110000000001011100000101001000100000000010100000101000010100110101000000000000000000010000000000100000001111000001101000001000000001000010000000000110000000010111010001011010010000000000000000000100000000110000001111000000000011111000000000000000000000010110100000001000110000000000000000000001100000100000000000001100000111010000010000111100100101110000001101011000000011111000111101100000010000100010000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000011110000001111100100100000000001010010000000110000000000001000001000011000000010000100000000000000101100011000010000000101010000000011010000100000111000110011000000001001010110010000001110100010100000000001000000000100001000110000101110101110100000000000101000000101000001100000000001000010100100100000100000000100000000010001011001000010010011000000001100000001100000000000010010001101001010010000001000000000010111000000000000010100000000001011000000110001100001100011000000001111000010000011000000001101000001000100000000000000110010100110001100000001100000000001010010000000000000000001000001100011111000010100001000000111100010000001000001010000100000000011100101001111010000001001000000000111010001100001001010101100000000000000010000000000001100110000000000000000011000110001100011000101000011000000000001001000011000001000000100110000000000000000000000000011011000000000000000000001000000101100000010010100000010011100000001000000101111111000011100010000000000000100000000100100000001000000000001010000000010000000000110111100100010000000000100101001111010001000000000100000000011010100000011100000000010100000011010000000100101110000000000000011000010001001001000001010000000001011011000000000100000110000110100011100100001110000100100100010101000000100000000010000000000000000000000000000000001000100001100100110011100000000000000010000000100000110000000000110000001000110000100000100000001100110001000000000001110010010000000001000010010111001100000100101111011000000011101000000011000000111100000000000101000110010000000001111011101001100000011100000000010100010000000000001110100000010000100000000000000000110010010001000001000000000011001000011100000100000010100000101100000000000000000101010000011000000000011000000000111001100000000000000010010111111110000000001011000000000000000000001000010000000000000000000000010000101000000010110010000000000000010101111110000001101000000111010000011100000000001100000000100001011000000110000000000000000000000000000010000000101000000000110000110010000001000000000111001000111000010000001110000000000000000100001010000000000000001010001100000000101111011100000000000100001110100000101110000010100000010111110010100000001101100001001110000000010000000000001010110000110001011010010000010010000000000000101001110000000000000000000000000000001010110001100110100011100100100000000110000000000101000001011010110000000000100011100001110100000010000110111111110000000010110000000000000000010000000001000000101010000100001000010001000100100000000010110110001111110100000000000000010000010110000100011010000001000000000010000001000110000011000100100100000001010101111000000000000000000000101100000001011000000000000000001010000001000010100000001000000000000001001110101110101000010100001001000010000000000010000000001000000000000000000000110100000111000000010101111000000100101111110101110110000000111010000000010000001010110000001100000000000010101010010000000011110100000000001000000000001101000100001000010010000001010100110101000001010111010000000001100110000000010000000000010100000000000010000000000010000000000000000000000000000000101100000001000100011100010001000011000100000000000010000111110000000111100000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000000100001101001100000111000000011000000000000000011100000000000000000001001001000000111101100001100000000100111011000000000000000111110110000000000100000000001100000010100010100000100000000000000000000011111100110100001000000000100011010000011100000000001001101111101100011010100000000100100011000000010010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000010100100010000001000000101000000000000000110010000000000111100000000000001100011100000010010011100010011010000000000000000000101001000000010110000010000100000000001000000000000000000010001000000000011",
	"0000001101000101101110100110000100101001110000100000010000001011111100001001000000000000110001000010110111000000011001101011011000000000100000000010110000010101000000100110110000111101000000010000000000000111111000000100000000011000000000000011000010000000000001011100000001000001011010110000001111100001010110010001110000000000010000001110101100000010000100000001010101000000001001000000001100000001101000100011111000001011011001110010010101000000000000000000110101110000000000000000010010110001000000001010110110110000100000000001100000001111100000001000010000100000100010000000010010000000000000000000000000000000000100111000010000000101000000000010010010010010010100000000000001100000000001100000000000000000100000000000010100111101001010000000000000000101100000000011011000000011011000011100001001101100000000000000000010101010101001001100011010000001000011000001010000010000000100010000001000000000001100000000010011010100000111100010010000001110010000000000100000010000000000100000000101100010001010101000010000010100100000100000100000000011110000000000000001000111110000110100000000000000000000011100000000001011010000010110000000000101101000000001000000000011111010000010100101110000011000000000101000000100001100000111000111000000010100000000000000001100100000000000100000101100001110101111100011100000000000100000000000000000000000001110000000001110000000000100000000000000010000000110000000000000000100001000000000000101011000000000000001010000000000100101000000110100000000001100101000000000111000101011000001101000000000111101100010000010000001000000000100011100000110110001111100000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000000000001010010000100110100000000000000000000011001100001100000000000000000000011000000000001100000000000010000000000110010000000000000100010000000000111000000000110000010000000011100001000000100000010000001010000001010110000011000110000000000001101010000000000000100110000000000100000001001000000000000100001011111011100000000000000010011000000000000010111000000100101000000000000000001100000000100000000100000000000110000001000101100111101100111100001011001100000000101101001110011001101000100010000000000000001100000011000100000100110000010000000100000000110000000100000000000000010000000100100100000000100000000000010100000001000000100010000000011000000000010000011001000101010100000010101101010000000000000000011100110001011110000001111001010101101000101000011111100000100010110100000000001101000000000000000001101000100000000000000000011100110110000000000001000000001011000100011100000010000000101000001011000000000000000011010011001011000010100101100000110000000000001000001000100000010000000000010100100100000011110001000000000000100011100111111000110000110010000001010000000000000000000011000100100100000011100010000000001100101001111010111000000000100000100000000101100001001111000000101011001010010100000000000000111100001011101100101100000010000000000111110000000000000001000001000100000000000000101000000010000000100001000000000010000000111000110110110111000000100011010100001000010110010000000001100000101000001000000100100000010000000011100000111001100000001110011000100000110000111100000011100001000001101010100000110000011111000000010110000000001010101010100000101000010001000100000001100000000001000000100000000000000010000001101100011001100001000000000000100000000011111100001010100001100000110001011101010111000000000000001100000100100100000000000001100001100000000000111100011000000101111010110000000010011000100000010000000000010000100000001000011000100000000000000000001001111010000000000001011101100100000001100000000010000001001000000100000000000000001110000000000000000010111000000001010000000111010001110110000000000011100100000000000010110000001000000000100010000000000000101100000000001011001101110110100000000000100000000000000011010001111111001101001011000001111001110000100001001100001001001101001000001100000000000000101001100010000110010000110001001100000001000101010000000000000000000111000111011100100100010000000010000000000001010111000010000101011100100000000000011000000000100100000001101110000000000011100000000010000000000000000101000001111000001100000001101101001001000100100001011010111101001000000110000100000000000011100101000000000000000100000000000000000000000000010001010100001001111100011000000111000000000010011000000000000000000000010000000000000000000000001110110100000000010000000010100000000000000000001111101100100000000000001000000010000001000000110010000000000000000000000110000000000000110001010010010000000001100000010101011110010101010100000000000001100000000000000001101101000001100000011010111011100111000010000001101011011000000010000000000000000000011000100000000000000000001000001100000100110110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000011000000000000010001110001110011000000010000000010100000000001000111111000000000000000000010000010100110110100000010100010011110000000100000100001000000000000100000000100000001110010011011100000000000100000000101000100010100010101010000000100110100011000000000000001001011100001111100001000010000000000001000000000010001010000000000010010110000000111001111101001101101011011000000000000111100000000010000000001011000000000001000100001100100000000011100001100000000011000000000001100010000010010000000011000000000100000000000010001011100000001101100011110111010011101000000100110100101000000100000010000000011110000101101101001100011100000000100001000000000010000000010010011010000000000110000000000000000001000000011011101000101100000000100100100010010000000000110010000101110000000110001011111101110000000001011100000101001000100000000010100000101000000100110101000000000000000000010000000000100000001111000001101000001000000001000000000000000010000000010111010001011010001000000000000000000100100000110000101111000000000011111000000000000000000000010110100000001000110000000000000000000001100000100000000000001100000111010000010000111101100101110000001101011000000011111000111101100000010000101000000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000011110000001111100100100000000001010010000000110000000000001100001000011000000010000100000000000000001100011010010100000101010000000011010000100000111000110011000000001001010110010000100110100010000000000001000000000100001000110000101110101110100000000000101000000101010001100000000001000010100100100000100000000000000000010000011001000010010011000000001100000001100000100000010010001101001010010000001000000000110111000000000000010000000000001010000000110001100001100011000000001111000010000011000000001101000001000100000000000000110010100110001100000001100000000001010010000000000000000001000001100011111000010100001000000111100010000001000001010000100000000011100101001111010000001001000000000111010001100001001010001100000000000000010000000000001100110000000000000000011000110001110010000101000011000000000001000000011000011000000100110000000000000000000000000011011000000000000000000001000000111100000010010100000010011100000001000000101111111000011100010000000000000100000000100100000001000000000001010000000010000000000110111100100010000000000100101001111010001000000000100000000011010100000011100000000010100000001010000000100101110000100000000011000000000001001000001010000000001011011000000000100000110000110101011100100001110000100100000010101000000100000000000000000000000000000000000000000000000100001100000110011100000000000010010000000100000110000001000110000001000110000000000100000001100110001000000000001110010010000000001000010010111001100000100101111011000000011101000000011000000111100000000000111000110010000100001111011101001100000011100000000011100010000000000001110000000010000100000000000000000110010010001000001000000000011001000011100000100000010100000101100000000000000000101010000011000000000011000000000111001100000000000000010010111111110000000001011000000000000000000001000010000000000000000000000010000100000000010110010000000000000010101111110000001101000000111010000011100000000001100000000100001011000000110000000000000000000000000000010000000101000000000110000110011000001000000000111001000111000010000001110000000000000000000001010000000000000001010001100000000101111011100000000000100001110100000101110000010100000010111110010100000001101100000001100000000010000000000001010110000110001011010110000010010000000000000101001110000000000000000000000000000001010110001100110100011100100100000000100000000000101000001011010110000000000100011100001110100000010000110011111110000000010110000000000000000010000000000000000101010000100001000010001000100100000010010110110001111110100000000000000010000010110000100011010000001000000000000000001000110000010000100100100000101010101111000000000000000000000101100000001011000000000000000001010000001000010100000001000000000000001001110101110101000010100001001010010000000000010000000001000000000000000000000110100000111000000010101011000000100101111110101110100000000111010000000010000001010110000001100000000000010101010010000000011110100000000001000100000001101000100001010000010000101010100110101000001010111010000000001100110000000010000010000010100000000000010000000000010000000000000000000000000000000101100000001000100011100010001000011000100000000000010000011110000000111110000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000100100001101001100000111000000011000000000000000011100000000000000000001001001000000111101100001100000000100111011000000000000000111110110000000000100000000001100000010100011100000100000000000000000000011111100110100001000000000100011010000011100000000001001101111101100011010100000000100100011000000010010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000010100100010000001000100101000000000000000110010000000000011100000000000001100010100000010110011110010011010000000000000000000101001000000010110000010000100000000000000000000000000000010001000000000011",
	"0000001101001101101110100110000100101001110000100000010000001011111100001001000000000100110001000010110111000000000001101011011000000000100000000010110000010101000000100110110000011111000000010000000000000111111000000100000000111000000000000011000010000000000101011100000001000001011010110000001111100001010111010001110000000000010000001110101100000010000100000001010101000000101001000000001100000001101000100011110000001011011001110010010101000000000100000000110101110000000000000000010000110001000000001010110110110000100000100001100000011111100000001000010000100000100010010000010010000000000000000000000000000000000100111000010000000101000000000010010010010010010100000000100001100000000001100000011000000000100001000000010100111100001010000000000000000101100000000011011000000011011000011100001001001100000000000000000010101010101001001000011000000001010011000001000000010000000100010000001000000000001100000000010011010100000111100010010000001110010000000000100000011000000000100000000101100010001011101000010000010100100000100000100000000011110000000000000001000111110000110100100000000000000000011100000000001011010000011110000000000101101000000001000000000011111010000010100101110000111000000000101000000100101100000111000111000000010000000001000000001100100000010100000000101100001110101111100011100000000000100000000000001000000000001110000000001110001100000110000000000000010000000110000000000000000100000000000000000101011000000000000001010000000000100101000000110100000000001100101000000000111000101011000001101000000000111100100010000010000001000000000100011000000110110001111100000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000000000001010010000100010100000000000000000000011001100001100000000000000000000011000000000001000000000000010000000000110010000000000000000010000000000111000000000110000010000000011100001000000100000010000011000000001010110000011000110000000000001101010000010000000100110000000000000000001001000000000000100001011111011100000000000000010011000000000000010111000000100101000000000000000001100000000100000000000000000100110000001000101100111101100111100001011001100000000101101001110111001101000100010000000000000001100000011000100000100110000010000000100000010110000000100000000000100010000010100100100000000100000000000010100000001000000100010000000011000000000110000011001000101010100000010101001010000001000000000011100110001011110000001111001010101101000101000011111100000100010110000000000001101000000000000000001101000100000000000000000011100110110000000000001000000001011000100011100000010000000101000001011000000000000000011010010001011000110100101100000110000000000001000001000100000010000000000010100100100000011110001000000000000100011100011111000110000110010000001010000000000000000000011000100000100000011100110000000001100101001111010111000000000000000100000000101100001011111000000100011000010010100000000000000111100001011101100101101000010000000000111110000000000000001000001000000000000000011101000001010000000100001000000000011000000110000100110110111000000100011010100001000010110010000000101100000101000001000000000000000010000001011100000101001100000001110011000100000110000111100000011100001000001101010100000110000011111000000010100000000001010101010100000100000010001000100000001100000000001000000000000000000000010000001101100011001100001000000000000100000000011111100001110110001100000110001011101010111000000000000011100001100110000000000000001100001100000000000111100011000000101111010110000000000011000100000010000000000010000100000001000011000000000010000000000001001111010000000000001011101100100000001100000000010000001000000000100000000000000001110000000010000000010111000000001010000000111010001110110000000000011100100000000000010110000001000000000100010000000000000101100000000001011001101110010100000000000100000100000001011010001111111001101001011000001111001110000100001001100001001001101001000011100000000000000101001000010000110010000110101001000000001000101010000001000000000000111000111010100100100000000000010000000000001010111000010000101011100100000000000011000000000100100000001101110000000000001100000000000000010000000000101000001011000001100000001101101001001000100100001001010111101001000000110000100000010000011100101000000000000000100000000000000000000000000010001011000001001111100011000000011000000000010011000000000000000000000010000000000010000000000001110110000000100010000000010100000000000000000001111101100100000000000001000000010000001000000110010000000000000000000000110000000001000110001010010010000000001100000110101011110010100010100000000001001100000000000000001101101000001100000111010111011100111000010000001101011011100000010000000000000000000011000100000000000000000001000001100000100010110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000011000000000000010001110001110010000000000000000010100000000001000111111000000000000000000010000010100110110100000010100010011110000000110000110001000000000010100000000100000001110010001011100000000000100000000101000100010100010101010000000100110100011000100000000001001011100001111100101000010000000000001000000000010001010000000000010010110000000111001111101001101101011011000000000000111100000000110000000011011000000000001000100001100100000000011100001100000010011000000000001110010000010010000010011000000000100000000000110001011100000001101100011110111010011101000000100110100101000000000001010000000001110000101101101001100111100000000100001000000000010000000010010011010000000001110000000000000000001000000011011100000101100000000100100100010010000000000110000000101110000000110001011111101110000000001011100000101001000100000000010100000101000010100110101000000000000000000010000000000000000001111000001101000000000000001000010000100000110000000010111010001011011000000000000100000100100100000110000101011000000000011111000000000000000000000010110100000001000110000000000000000000001100000100000000000001100000111010000010000111100100101110000001101011000000011111000111101100000010000101010000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000011110000000111100100100000000001010010000000110000001000001000001000011000000010000100000000000000101100011000000000000101010000000011010000100000111000110011000000001001010110011000101110100010000000000001000000000100001000110000101110101110100000000000001000000101000001100000000001100010100100100000110000000100000000010000011001000010010011000000001100000001100000000000010010001101001010010000001000000000010111000000100000010100000000001010000000110001100001100011000000001111000010000011000000001101000001000100000000000000110010100010001100000001100000000001010000000000000000000001000001100011111000010100001000000111100000000001000001010000100000000011100101001111010000001001000000000111000001100001001010001100000000000000000000000000001100010000000000000000011000110011100000000101000011000000000001001000011000001000000100110000000000000000000000000011011000000000000000000001000000111100000010010100000010011100000001000001101111111000011100010000000000000100000000100100000001000000000001010000000010000000000110111100000010000000000100101000111010001000000000100000000011010100000011100000000010000000001010000000100000110000100000000011000010000000001000001010000010000011010000000000100000100000110100011100100001110000100100100010101000000100000000010000000000000000000000000000000001100000001100000110011100000000000010010000000100000110000001000110000001000110000000000100000000100110001000000000001110010000000000001000010010111001100000100101111011000000011101000000011000000111100000000000110000110010000100001111011001001100000011000000000011100000000000000000110000010010000100000000000000000110010010000000001000000000011001000011100000100000010100000101100000000000000000101010000011000000000011000000000111001100000000000000010010111111110000000001011000000000000000000001000010000000000000000000000010000101000000010110010000000000000010101111110000001101000000111010000011100000000001100000000100001011000000110000000000000000000000000000010000000101000000000110000110010000001000000000111001000111000010000001110000000000000000100001010000000000000000011001100000000101111011100000000000100001110100000101110000010110000010111110010100000001101100001001100000000000000000000001010110000110001011010010000010010000000000000101001110000000000000000000000000000001010110001100110100011100100100000000110000000000101000011011010110000000000100011100001110100000010000110111111110000000010110000000000000000010000000000000000101010000100001000010001000100100000010010110110001111110100000000000000010000010100000100011010000001000000000000000001000110000000000100100100000001010101111000000000000000100000101100000001011000000000000000001010001001001010100000001000000000000001001110101110101000010100001001000010000000000010000000001001000000000000000000110100000111000000110101111000000100101111110101110100000000111010000001000000001010110000001100000000000010101010010000000011110100000000001000000000001101000100001010000010000101010100110101000001010111010000000001100010000000010000010000010100000000000010000000000010000000000000000000000000000000101100000001000100011100010001000011000100000000000010000111110000000111100000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000100100001101001100000111000000011000000000000000011100000000001000000001001001000000111101100001100000000100111011000000000000001111110110000000000100000000001100000010100011100000100000000000000000000011111100110100001000000000100011000000011100000000001000101111101100011010100000000100100011000000010010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000000100100010000001000000101000000000000000110010000000000111100000000000001100011100000010100011110010011010000000000000000000101001000000010110000010000100000000000000000000000000000010001000000000011",
	"0000001101000101101110100110000100101001110000100000010000001011111100011001000000000100110001000010110111000000010001101011011000000000100000000010110000010101000000100110110000011111000000010000000000000111111000000100000000111000000000000011000010000000000001011100000001000001011010110000001111100001010110010001110000000000010000001110101100000010000100000001010101000000101001000000001100000001101000100011111000001011011001110010010101000000000100000000110101110000000000000000010100110001000000001010110110110000100000000001100000001111100000001000010000100000100010010000010010000000000000000000000000000000000100111000010000000101000000000010010000010010010100000000100001100000000001100000001000000000100001000000010100111100001010000000000000000101100000000011011000000011011000011100001001101100000000000000000010101010101001001100011010000001010011000001000000010000000100010000001000000000001100000000010011010100000111100010010000001110010000000000100000010000000000100000000101100010001000101000010000010100100000100000100000000011110000000000000001000111110000110100100000000000000000011100000000001011010000011110000000000101101000000001000000000011111010000010100101110000110000000000101000000100001100000111000111000000010000000000000000001100100000000100000000101100001110101111100011100000000000100000000000001000000000001110000000001110000000000110000000000000010000000110000000000000000100000000000000000101011000000000000001010000000000100101000000110100000000001100101000000000111000101011000001101000000000111100100010000010000001000000000100011100000110110001111100000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000000000001010010000100010100000000000000000000011001100001100000000000000000000011000000000001000000000000010000000000110010000000000000100010000000000111000000000110000010000000011100000000000100000010000011010000001010110000011000110000000000001101010000010000000100110000000000100000001001000000000000100001011111011100000000000000010011000000000000010111000000100101000000000000000001100000000100000000000000000000110100001000101100111101100111100001011001100000000101101001110111001101000100010000000000000001100000011000100000100110000010000000100000010100000000110000000000100010000010100100100000000100000000000010100000001000000100010000000011000000000110000011001000101010100000010101001010000000000000000011100110001011110000001111001010101101000101000011111100000100010110000000000001101000000000000000001101000100000000000000000011100110110000000000001000000001011000100011100000010000000101000001011000000000000000011010010001011000010100101100000110000000000001000001000100000010000000000010100000100000011110001000000000000100011100011111000110000110010000001010000000000000000000011000100100100000011100110000000001100101001111010111000000000000000100000000101100001011111000000000011001010010100000000000000111100001011101100101100000010000000000111110000000000000001000001000000000000000000101000001010000000100001000000000011000000111000110110110111000000100011010100001000010110010000000001100000101000001000000000000000010000000011100000101001100000001110011000100000110000111100000011100001000001101010100000110000011111000000010110000000001010101010100000101000010001000100000001100000000001000000100000000000000010000001101100011001100001000000000000100000010011111100001110110001100000110001011101010111000000000000001100000100100000000000000001100001100000000000111100011000000101111010110000000010011000100000010000000000010000100000001000011000000000000000000000001001111010000000000000011101100100000001100000000010000001000000000100000000000000001110000000000000000010111000000001010000000111010001110110000000000011100100000000000010110000001000000000100010000000000000101100000000001011001101110010100000000000100000000000001011010001111111001101001011000001111001110000100001001100001001001101001000011100000000000000101001000010000110010000110101001000000001000101010000000000000000000111000111010100100100010000000010000000000001010111000010000101011100100000000000011000000000100101000001101110000000000011100000000010000000000000000101000001111000001100000001101101001001000100100001011010111101001000000110000100000000000011100101000000000000000000000000000000000000000000010001010100001001111100011000000011000000000010011000000000000000000000010000000000000000000000001110110000000000010000000010100000000000000000001111101100100000000000001000000010000001000000110010000000000000000000000110000000001000110001010010010000000001100000010101011110010101010100000000001001100000000000000001101101000001100000011010111011100111000010000001101011011000000010000000000000000000011000100000000000000000001000001100000100110110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000011000000000000010001110001110010000000000000000010100000000001000111111000000000000000000010000010100110110100000010100010011110000000110000100001000000000000100000000100000001110010001011100000000000100000000101000000010100010101010000000100110100011000100000000001001011100001111100001000010000000000001000000000010001010000000000010010110000000111001111101001101101011011000000000000111100000000110000000001011000000000001000100001100100000000011100001100000010011000000000001110010000010010000010011000000010100000000000010001011100000001101100011110111010011100000000100110100101000000000001010000000001110000101101101001100011100000000100001000000000010000000010010011010000000000110000000000000000001000000011011100000101100000000100100100010010000000000110000000101110000000110000011111101110000000001011100000101001000100000000010100000101000010100110101000000000000000000010000000000100000001111000001101000000100000001000010000100000110000000010111010001011011001000000000000000100100100000110000101011000000000011111000000000000000000000010110100000001000110000000000000000000001110000100000000000001100000111010000110000111101100101110000001101011000000011111000111101100100010000101010000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000011110000001111100100100000000001010010000000110000000000001000001000011000000010000100000000000000001100011000010100000101010000000011010000100000111000110011000000001001010110010000101110100010000000000001000000000100001000110000101110101110100000000000101000000101000001100000000001100010100100100000100000000000000000010000011001000010010011000000001100000001100000100000010010001101001010010000001000000000010111000000000000010000000000001010000100110001100001100011000000001111000010000011000000001101000001000100000000000000110010100010001100000001100000000001010010000000000000000001000001100011111000010100001000000111100000000001000001010000100000000011100101001111010000001001000000000111010001100001001010001100000000000000000000000000001100010000000000000000011000110001100000000101000011000000000001001000011000001000000100110000000000000000000000000011011000000000000000000001000000111100000010010100000010011100000001000001101111111000011100010000000000000100000000100100000001000000000001010000000010000000000110111100100010000000000100101001111010001000000000100000000011010100000011100000000010000000001010000000100000110000100000000011000010000000001000001010000010000011010000000000100000110000110101011100100001110000100100100010101000000100000000010000000000000000000000000000000001100000001100000110011100000000000010010000000100000110000001000110000001000110000000000100000000100110001000000000001110010010000000001000010010111001100000100101111011000000011101000001011000000111100000000000111000110010000100001111011101001100000011000000000011100000000000000000110000010010000100000000000000000110010010001000001000000000011001000011100000100000010100000101100000000000000000101010000011000000000011000000000111001100000000000000010010111111110000000001011000000000000000000001000010000000000000000000000010000101000000010110010000000000000010101111110000001101000000111010000011100000000001100000000100001011000000111000000000000000000000000000010000000101000000000110000110010000000000000000111001000111000010000001110000000000000000100001010000000000000001011001100000000101111011100000000000100001110100000101110000010110000010111110010100000001101100001001100000000000000000000001010110000110001011010010000010010000000000000101001110000000000000000000000000000001010110001100110100011100100100000000100000000000101000011011010110000000000100011100001110100000010000110011111110000000010110000000000000000010000000000000000101010000100001000010001000100100000010010110110001111110101000000000000010000010110000100011010000001000000000000000001000110000010000100100100000001010101111000000000000000100000101100000001011000000000000000001010001001001010100000001000000000000001001110101110101000010100001000010010000000000010000000001001000000000000000000110100000111000000010101111000000100101111110101110100000000111010000001010000001010110000001100000000000010101010010000000001110100000000001000000000001101000100001010000010000101010100110101000001010111010000000001100110000000000000010000010100000000000010000000000010000000000000000000000000000000101100000001000100011100010001000011000000000000000010000111110000000111110000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000100100001101001100000111000000011000000000000000011100000000001000000001001001000000111101100001100000000000111011000000000000001111110110000000000100000000001100000010100011100000100000000000000000000011111100110100001000000000100011000000011100000000001000101111101100011010100000000100100011000000010010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000000100100010000001000000101000000000000000110010000000000111100000000000001100011100000010100011110010011010000000000000000000101001000000010110000010000100000000000000000000000000000010001000000000011"
	); --six test class HVs, one for each vowel
  	variable test : testarray := ("0000001101001101101110100101000100001001100000100000000001001011111100001001000000000000110001000010110111000000010001101011011000000000100000000010110000010101010000100110110000011111000000010000000000000011111010100100000000111000000100000011000010000000000001011100000001001011001010110000001111100001100111010000110000000000010000001110101000000010000000100000010101000000101001000000001100000000101000000011110000001011001001110010010101000000000100001000110001110000000100000000010000100001000000001110110110110000100000100001100000001011100000001000010000000000100010010000010010000000000000000000000000000000000100111000010000000101000000001010010001010001010100000000100001100000000001100000001000000100100001000000000100111100001010000000000000000100110000000011011000000011011000010100001001101100000000000000000010101010000001001100011010000001010011100001100000000100000100010000001000000000001001000000010111011000000011100010000000011110000000000100000100001000000001100000000101100010001001101000010000010100100000110100101000000010110000000000000001000011110000110100100000000100000001011100000000000011010000011110000000000101101000000001010000000011111010000010100101110000101000000000101000000100100100000111000111010000001000000001000000101000100000010100000000100101001110101111100011100000000000100000000000001000000000001110000001001111001100000010000000000000010000000100001010000100000100000000000000000101011000000000000001010000010010100101000000110100000000001100101000000010111000111011000001101000000000111100100010000010100000000000010000011100000111010001111100000000000001000000001100010010000000000000011100000000000000000001100000000000000001000000000101000001010010000100010100000000000000000000011001110001100000000000000000000010000001100101000000000000010000000000110010000000010000000010000000000111000000000110000010000000111100000000000100000110000011000000000010101000010000100000000000000101010000010000000100110000000000000000001001000000000001010001011111011100000000000000010001000000000000000111000000100101000000000000000101100000000100000000000000000000110100001000111100111101100111000001011001100100000111101001110100001101000100010000000000000001000000011000100000000100000010000000100000011110000000110000000000100010000010100100100000000000000000000010100000001000000000010000000011000000000110000011001100101010100000010101001010100010000000000001110000001011110000101111001010101101000101000011111100000100010111000000000001001000000000001000001101000000100000000000000111100110110000000000001000000001011000100011100010100000001101000001011010000001000000011010010101011000010100101100000110000000000001000001000100000010000000000010100000100000011110001000000000001100011100011110000110000110010001011010100000000000000000011000100000100000010100110000000001100101001111010111000000000000000100000000001100000011111000010000011000010010100000001001000111100000011101100101100100010000000000111110000000000000011000000000000000000000010101000001000000001100001000000000011000000010000100110110111000000100011010100001000010110010000000101100000101100001000000000100000010000001011100010100001100000001111011100100000110010111100000011100001100001101010100000110000111111000000010110000000001010101010100000101000000001000100000001100000000001100000010000000000000010000001101100011001100001000000000000100000010011111100001110010001010010110001011101010011000000000000001100000101100000000000000001100001100000001000101100011000000101111010110000000010011000100000010000000000010000100000011000011000000000000000000000001001111010000000000001011101100000000001100000000010100001000000000100000000010000000100000000000000000010111000000001011000000111000001110110000000000011100100000001000110110000001000000000100010000000000000101100000000001010000100110010100000000000000000000000000111010001110011001101000000000001110001110000100001001000001001001101001010011100000000000000101001100010000110010000110101001000000001000101010000001001000000000111000111010100100100010000000010010001000010010111000010000101011100100000000110010000000000000100001001101110000000100011100000000000000000000010000101000001111100001100000001101100001011000100000001011010111101001000000100000110000011000110100101000000000000000000000000000000000000000000000001001100000001111100000000000111000000000010011100000000000000000000010000000000010000000000001110110000000000010000000010100000000000000000001111100100100000000000001000000010000000000000110010001000000000000010000110000000001000110001010010010000000001100000000000011100010100010100100000001001100000000000000001101101010001000001011010111010100111000010000001101011010000000010000010000000000000011100101001000000000000010000001100000000110110101010000000000000001100000000000000101000000000000001000001110000001100010000000000000000000001010000000000011000000000000000001110001110010000000000000000010100000000001000011110000000000000000001010000010100110110110000110100010011110000000110000000001000000010010100000000100000001010010101011100000000001100000000111000100010100010100010000000100110100010100100000000001001011100001111100000001000000000000000000000000000001110000000000010010110000000111001111101001101101011011000000000000110000100000110000000001011000000000001000100001100100000001010100001100000011011000000000001010010000000010000000011000001010000000000000010001011100010001101100011110111010010101000010100110100101000000001001010001000101110000101101101001100011100000001110101000000000000000000000010011010000000001110000000000000010001000000011011100000101100000000000100000000010000000000110000000101100000000110110011011101110000000001011100000101001000100000000110100000001000010100110101000000000000000000011000000000000000001111000001101000001000000001000010000100000110000001010111010001011001000000000000100000100100100000110000101011000000010011111000010000000000000010000110100000001000010000110000000000000011110100000000000000001010000111010010110000101100100100100000001101011000000011111000111101100100010000011011000101010001011000000110000001000001010011001110110000000000000111000100100101100110000000011110000000111100100100100000001010010000100110000001000001000000000011000000010000100001000000100001100011000000100000101010000000011010000100001111000110010000000001001010111011000100110100110000010000001000000000100000000111000101110101110000100000101001000000101000001100000000001100010100100101000110000010100000000010000011001000010010011000000001100000001100000100100010010000101001010010000001000000001010111000000100000010000000000001010000100110001100001100011001000001111000001000011000000001101000001010100000000000000110010100010001100000001100100000011010000000000000000000001000001110001110000010100000000000111100000000001000001010010100000000011100101001111000000000001000000000111010001100001001010001000000000000000100000000000000101010000000000000000011000010001100000000001000011000000000001001000011000001000000000110000000000000000000000000011011000000000000000000001000000111100000011000100000010011100000000000000101111111000011100000000000000010100000010100100000001000000000001010000000001000000000110111100000010000000000100101000110010001000000000100010000011010100000011100000000010000000001010000000100000111000100000000011000010001000001000000010000010000011010000000100100000100000110101011000000011110000100100000010101000000100000000010000000000000000000000000000000001100001001000100110011100000000000010010010000100000100000001000100000001000110000010000100000000100100001000000000001110010000001000001000010010111001100000100101111011000000111101000001011000000101100000000000110000010010000100001111011001001100000011000000000011100001000000010000100100010010000100000000000000000110010010000000001000000000011001000011100010100000010100000101010000000000000000100000000011000000000011000000000101001100000000000000010010111111110000000001011000000000000000010011000010000000000000000000000010000001000010010110010000001000000010101111010000001101000100111010000011100000000001100000000000001011000000111000000000010000000000000100010000000101000000000110000110010000001000000000111001000111000010000001110000000000000000100001000000000000000011011000100000000101111011100000000010100001110100000001110000010010000010111100010100000000101100001010100000000101000000000001010111000110011011010000000010010000000000000101000110000000001000000000000010000001010110001100110100001100100100000000100000000000101000011011010110000000000100011100001110100000010000110111111110000000010110000000010000001010000000011000000001010010100000001011010000100000010010010110110001111110101000000000000010000010101001000011000000001000100000000000000000110000000000100100101000001010101111000000000000000100000101100000000001000000100000000001000001001001010100000000000000000000011001110101110000000010100001000010010000000000010000000001001100000000000000000110000010011000000110100111000000100101111100101110100000000011010000001000000001000110000001100000000000010101010000000000001110100000000001000000000001101010100001000000010000100010100110100000001010111010000000001100000000000000000010000000100000000000010101000100010000000000000000000000000000000010100000001000000011100010001000011000000000000001000000011110000000111110000001110101100000000100000001110110000111100100000000000001000001100010000000000000011010000100010101101001100000111000001011000000000000000011100000000001000000001001001000000111101000001100100000100111011000000000000001111110110000000000101000000001100000000101011100000100000000000000100000011111110010100011000010000100011000000011100000000001000101111100100011010100000000100100011000000010000110111110110110000000111000110110000000000000000000100000000000100100010010100011010010001010000000100100010000001001000101000000000000001110010000000000111100000000000001100001100000010100111110110011010000000000000000000101001000000010010010010000100000000000000000000000000000000001000000000001",
	"0000001100000101101110100110000100101001110000100000000000001011111100011001000000000100110001000010110111000000010001101011011010000000100000000010110000010101010000100110110000011111000000010000000000000111111010000100000000011000000000000011011010000000000001011100000001000001011010110000001111100001010110010000110000000000010000001110101100000010000100100001010101000000101001000000001000000001101000100011111000001011011001110010010101000000000100000000110001110000000000000000010100110001000000001010110110110000100000000001100000001011100000001001000000000000100010010000010010000000000000000000000000000000000100111000010000000101000000000010010101010011010100000000100001100000000001100000001000000000101001000000000100111110001010000000000000000101100000000011010000000011011000010100001001101100000000000000000010101010101001001100011010000001010011100001100000010000000100010000001000000000000000000000010011011000000011100010010000001110000000000000100000010000000000100000000001100010001001101000010000010100100000100000100000000011110000000000000001000011110000110100100000000000000000011100000000000001010000011110000000000101101000000001010000000011111010000010100101110000110000000000101000000100000100000111000111010000011000000000000000001100100000000100000000101100000110101111100011100000000000000000000000001000000000001110000100001111000000000010000000000000010000000110000000000000000100000100000000000101011000000000000000010000000010100101000000110100000000001100101000000000111000101011000001101000000000111100100010000010100001000000000000011100000110010000111100000000000001000000001100010010000000000000011100000000000000000001100000000000000001000000000001000001010010000100010100000000000000000000011001100001100000000000000000000011000000000101100000000000010000000000110010000000000000100010000000000111000000000110000010000000011100000000000100000010000011010000001010110000011000110000000000001101010000000000000100110000000000100000001001000000000000110001011111011100000000001000010011000000000000010111000000100101000000000000000101100000000100000001000000010000110100001000101100111101100111100001011001100100000111101001110111001101100100010000000000000001100000011000100000000110000010000000100000010100000000110000000000100010000010100100100000000100000000000010100000001000000000010000000011000000000110000011001100101010100000010101101010000000000000000001110110001011110000001111001010101101000101000011111100001100010110100000000001101000000000000000001101000100000000000000000011100110110000000000001000000001011000100011100000110000001101000001011000000001000000011010010001011000010100101100000110000000000001000001000100000010000000000010100000100001011110001000000000000100011100011111000110000110000000011010000000000000000000011000100100100000011100110000000001100101001111010111000000000000000100000000001100001011111000000000011001010010100000000000000111100001011101100101100100010000000000111110000000000000001000000000000000000000000101000001010000000100001000000000011000000111000110100111111000000110011010110001000010110010000000001100000101100001000000000100000010000000011100010111001101000001111011100100000110010111100000001100001100001101010100000110000011111000000010110000000001010101010100000101000010001000100000001100000000000000000110000000000000010000001101100011001100001000000000000100000010011111100001100010001010000100001011101010011000000000000001100000110100000000000000001100001100000000000111100011000000101111010110000000010011000100000010000000000010000100000001000011000000000000000000000001001111010000000000000001101100000000001100000000010000011001000000100000000000000000110000000000000000010111000000001010000000111010001110110000000000111100100000000000010110000001000000000100010000000000000101100000000001011001101110010100000000000100001000000001011010001111111100101001011000001111001110000100000001110001000001101001010011100000000000000101001000010000110010000110101001000000001100101010000000100000000000111000111010100100100001000000010000000000001010111000010000101011100100000000010011000000000000101001001101110000000000011100000000110000000000010000101000001111100001100000001101101001001000100100001011010111101001000000110000100000000000011100101000000000000000000000000000000000000000000010001001100001001111100010000000111000000000010011000000000000000000000010000000000000000000000001110110000000000010000000010100000000000000000001111101100100000000000001000000010000001000000110010100000000000000000000110000000001000110001010010010000000001100000010101011110010100010100100001001001100000000000000001101101000001000000011010111011100111000010000001101011011000000010000010000000000000011000101001000000000000010000001100000100110110101010000000000000001100000000000000101001000000000001000000110000001100010100000000000000000001010000000000000000000000000000001100001110011000000010000000010100000000001000111111000000000000000000010100010100110110110000110100010011110000000110000100001000000000000100000000100000001110010101011100000000000100000000101000000010100010101010000000100110100001000100000000001001011100000111100000000010000000000000000100000000001010000000000010010110000000111001111101001101101011011000000000000111100100000110000000001011000000000001000000001100100000000011100001100000010011000000000001110010000010010000000011000000010100000000000010001011100000001101100011110111010010100000000100110100101000000011001010000000001110000101101101001100011100000000110101000000000000000000000010011010000000000110000000000000000000000000011011101000101100000000000100100000010000000000110000000101110000000110010011111101110000000001011100000101001000100000000010100000001000000100110101000000000000000000011000000000100000001111100001101000001100000001000010000100000110000000010111010001011001010000000000000000100100100010110000101011000000010011111000010000000000000000010110100000001000110000000000000000000001110100000000000000001100000111010000110000111101100100100000001101011000000011111000111101100100010000001000000001010101011000000010000001000001010011001110110000000000000111000000100101000110000000001110000000111100100000000000001010010000100110000000000001100001000011000000010000100001000000000001101011010010100000101010000000011010000100000111000110011000000001001010111010000000110100110000000000001000000000100001000110000101110101110100000000000101000000101000001100000000001100010100100001000100000000000000000010000111001000010010011000000001100000000100000100100010010001101001010010000001000000000010111000000000000010000000000001000000100110001100001100011001000001111000011000011000000001101000001010100000000000000110010100010001100000001100100000001010010000000000000000001000000100011111000010100001000000111100000000001000001010000100000000011100101001111000000001001000000000111010001100001001010000100000000000000100000000000001100010000000000000000010000110001100100100001000011000000000001001000011000001000000000110000000000000000000000000011011000000000000000000001000000111100000010000100000010011100000000000001101111111000011100000000000000000100000000100100000001000000000001010000000011000000000110111100100010000000000100101001111010001100000000000000000011010000000111100000000010100000001010000000100010111000100000000001000010000000001000000010000010000011010000000000000000110000110101011100100001110000100100000010101000000100000000010000000000000001000000000000000000100000001100000110011100000000000010000000000100000110000001000110000001100110000000000100000000100110001000000000001110010000000000001000010010111001100000000101101011000000111101000001001000000101100000000000111000010010000100001111011001001100000011000000000011100011000000000000110000010010000100000000000000000110010010001000001000000000011001000011100010100000010100000001100000000000000000101010000011000000000011000000000111001100000000000000010010111111111000000000011000000000000000000011000010000000000000000000000010000001000000010110010000001000000010101101010000001101000000111010000011100000000001100000000000001011000000111000000000000000000000000000010000000101000000000110000110010000000000000000111001000111010010000001110000000000000000100001010000000000000011011001100000000101111011100000000000100001110100000000110000010110000010111110010100000000101100001001100000000100000000000001000111000110001011010010000010010100000000000101001110000000001000000000000010000001010110001100110100011100000100000000100000000000101000010011010110000001000100011100001110100000010000110111111110000000000110000000010000001010000000000000000101010000100001001010010000100100000010010110110001111110101000000000000000000010111001000011010000001000000000000000100000110000001000100100101000001010101111000000000000000100000101100000000011000000000000000001010001001001010100000001000000000000001001110101110101000010100001000110010000000000010000000001001000000000000000000110100010111000000010100110100000100101111110101110100000000111010000001100000001010110000001100000000000010001010010000000001100100000000001000000000001101010000001010000010000101010100110100000001010011010000000001100110000000000000010000000100000000000010000000000010000000000000000000000000000000100100000001000100011100010001000011000000000000000000000011000000000111110000001110101100000000000000001110110010111100100000000000000000001100000000000000000001010000100110101101001100000111000001011000000000000000011100000000001000000001001001000000111101100001100000000100011011000000010000001111110110000000000101000000001100000010101011100000100000000000000100000011111100010100010000000001100011010000010100000000001010101111101100011010100000000100100011000000001010110111110100110000000111001110111000000000100000000100000000000100100010010100011010011001010000000100100010000001001000001000000000000000110010000000000111100000000000001100001100000010110111110010011010000000000000000000101001000000000010000010000000000000000100000000000000000010001010000000001",
	"0000001101001101101010100010000100001001000000100000010000000011111100011001000000000100100001000010100110000000000001101011011000000000100000000010110000000101000000100110110000111110000000010000000000000111111000100100000001111000000000000010000010000000000101011000000001001000011010110000001111100001000111000001110000000000010000011100101100000010000110000001010101000000111001000000001100000001101000100011100001001011001001110010010101000000000100001000110001110000000100000000011000100001000000001110110110110000100001100001100000011111100010011000110000000000100010010000010010000000000000000000000000000000000000111000110000000101000000101010010000010000010100001000100001000000000001100000011000000000100001000100010100111000001010000010000000000101100000000010010000000010011000011100001001001100001000000000001010101010001001001000011000000001010011000001000000010000000100010010001000000000001010000000010001011100000111100010000000011110000000000000000000011000000000100000000101100010001001101000011000000100100000100000100000000000110000000000000000000111100000110100100000010100000000010100000000101011010000011000000000000100100000000001000000000111111010001010100101110000111000000001101000000000101100000111000111000000010000000001000000001000100000010100000000101100001110001111100011100000000000100000000100001000000000001110000011001110001100000110000000000000010000000110010100001000000100000000000000010001011000000000000000010000010000100101000000110100000000001100100000000000111000101011000001101000000010111100100010000010100000000010000100011000000110110011111100000000000000000000011100010010000000000000011100000000010001000001100000000000000001000000000000000001010010000100110100000000000000000000011001100101100000000000000000000010000001100101000000000000010000000000110010010000000000000010000000000111000000000110000010000000011100000100010100000110000011000000001010010001001000110000000001001101010000010000000100110000000000000000001001000100000000110001011111011000000000000000010010000000000000010111000000100101000000000000000001100000000000000000000000010100110000001000001100111101100110000101011001100000000101101000110011001101010100010001010000000000100000011000000000100110000010000000100000010110000000100000000000100010000010100100100000100000000000000110100000001000000100010000000011000010000110000011001000101010100000010101001010000001100000000010100011001011110001101111000010101101000100000011111110000100010100000000000000100000000000000000001101000100100000000011000011100110100000000000001100000001010000100011000010000000000100000001011000000000000000011010011000011000110100101100010110000011000001000101000100000010000000000010100000100000001110001000000000011100011000011110000110000110010001001010000001000000000000011000100000100000011100110001000001100101001111010111000000000000000101000000100100000011111000010100011000010000000000100000000111100001011101100101101000010000000000111111000000000000111000001000000000000000011001000001010000010100001000000000010100000100000100110110000000000100011010000001010010110010000000101100000101000000000000010000000010000001011100000001001000000001110011000100000100000111100000011100001000001101010100000110000111111000000010100000000000010101010100000100000010001000100000001100000000101000000000000000000010010001001101100011001100001000000000000100000000011111100001100100001000010110001011101010011000001000000011100001100010000000010000001100001000000001000111100011000000101111010110000010000011000100000110000000000100000100000000000011000000011010000000000001001111010010000000001011100100100000001100000000000110001000000000100000000000000001110000000010000000010000000000001010000100111001001110110000000010011100100010000000110110000000000000000100010000000000000101100000000001001001100110010100000000100100000100100001011000001110011001101001000000101000001110000100011001000001001011101000000111100000000000000101000000010000110010000110101001000000000000101010000001001000000000111000111000101100100000000001010000000000101010111100010000101011100100000000010011000000000100100000001101110000000100001100000000000000010000100000000000001001000101100000001101100101001010000100001000010111100001000000100000100001011000101100100000000000000000100000000000000000100000000010001011000001001111100001000000011000000000010011000000010000000001000010000000000010000001000011100110000000100010000000010100000000000000000001111100100100000000000001000000010000001000000110010000000000000000110000100000000001000110001010010010000000001100000010100011100010100010100000000001001100000000000000001101101110001100011111010111000100111000010000001101011011100000010000000000000000000011000100000000000000000001000001100000100000110101010000000000000011100000000000000101000100000000001000001110000001100000100000000000000000001010000000000011000000000000010001100001110010000000000000000010100000000001000111100000000001000000000010000010100110110100000000100010011110000000110000010001000100010010100000010100000000010010001010000000000000100000000101000101010100000101010000000000110100101000100000000001001011100001111000100100010000000000001000000000011001110100000000010010110000000111001111101000101101001011000000000000101100000000110000000011011000000000101000000001100100000010001100001100000010010000010000000010110000010000000010011000100000100000000000110001011100000001101100011110111010011100000000000110100101000000000001010000000001110000101101001001100111100000000110001000000000010000000010000011010000000001110000000000000000001000000011011100000111100000000100100000010000000000000110000000101110000000100101010011101110000000001011100010101001000000000001110100000101000010100000101000000000000000000010000000000000000001110000001101000000000000001000010000000000110000001010111110001010011000000000000100010100100000000110000001010000000000010111000000000000000000000000100000000001000010000000000000000000000100000100000000000001100000111010001010010011100000101110000001101011000000011111000111101100000010000111011001001010001011000000110000001000001010001000110110000000000000111000000100101000100000110011110000000111100100000000000001010010000000110000001000001000001000011000000010000100000000000100101100011000000000000101010000001011010000100000111000110001000000001001010110011000101110100000000100000001000000000100001000110000100110101110100000000100001000000100000001100000000001100010100100101010110000000100000000010000011001000010010011000000001100000001100001000000010010001101001010010000001000001000010111000100100000010100000000001011000000110001100000100011000000001111000010000011000000001101000011010100000010000000110010100010001100000111100000000011010000000000001100000001000001110001110000010100001000000111000000000001000001010010100000000011100101001110010000001001000000000111000001100001001010001100010000000000000000100000001100010000000000000000011000110011010000000001000011000000000001001000011000001000000100010000000000000000000000000011011000000000001100001101000000101100000011010000000010011100000001000001101000011000011100000000000000000100010000100000001001000000000001010000000000000000000110111100000010000000000100101000111010000000000000100010000011010100000011100000000010000000011010000000100000110000000000000011000010000001001000011010000010000001010000100000100000000000110100010000000001110000100000100010101000000100000100010000000000000000000000000000000011100011000000000110011100000000100010010010000110000100000000000100000001100110000100000100000000100110001000000000001100010000000000001000010000111001100000000001111011000000011101000000011000000111000000000000100000110010000100001111011000001100000010000000000010000000000010000001000100110000000100000000010000000110010000000000001100000000010001000011100000100000010100000100110000000000000000101010000001000000000011000000000011001100000000000000010010111111110000000001011000100001000000000000000010000000000000000000000010000100000000000110010000000000000010101111110000001101000100111010000011100000000001100000000100001011000000110000000000000010000000000000010000000100000000000010000110010000000000000000111001000111000010000001110100000001001000100001000000000000000000010001100000000101111011100000000000100001110000000100100000000110000010111000010100000001101100001111110000000010000000000001010110000110011001010010000010010000000000000101001110000000000000000000000000000001010110001100110100011100100100000000110000000000101000011011010110000000000000011000001110000000010000110101101110000000010110000000000000000010000000000000000101010000100001010010001000100100010010010110110001111110100000000000000010000010100001100011010000001000000000000000101000110000000000100100000000000010101111000000000000000100000101100000001011000000000000000001000001001001010100000000000000000000111001110101110000000010100001001000010000000010010000000001001000000000000000000110000000111000000110101111000000100101111000101110110000000111010000000010000001010111000001100000000000110101010000000000001110100000000001000000000001101000100001000000010000000110100110101000001010111010000000001100000000000010000000000010000000000000010000000001010000001010000000000000000000000101000000001000100011100010001001001000100000000001010000111110000000111100000001110001100000000100001001110110010111100100000000000000000001000000000000000000111010000000111001101001100001111000000011000000000000000001100000000001000000001001001000010111001000000100110000000111011000000000000110111110110000000000100000000001100000010100011101011100000000000000000000011111110110000010000010000100011000000011100000000001000100111100100011010100000000100100011000000010010110111110100110000000111001110110000000000100000000100000000000100100010010100011010001001010000000100100010000001000000101000000000000001110000000000000111100000000000001100011100000010000011110010011010000000001000000000101000000001110100000010000100000001000100000000000000000010001000000100011",
	"0000001101001101101010100101000100001001000000100000010000001011111100001001000001000000110001000010110111000000000001101011011000000000100000000010110000010101000000100110110000011111000000010001000000000011111000100100000000111000000100000011000010000000000101011100000001001011001010110000001111100001000111010001110000000000010010001110101000000010000000000001010101000001111001000000000100010000101000000011010000001011001001110010010101000000100100001000110001110000000100010000010000100001000000001110110110100000100001100001100000011111100000001000010000100000100010010000010000000000000000000000000000000000000100111000010000000101000000000010010000010000010100001000100001100000000001100000011000000000100011000100010100111100001010000000000000000100110000000011011000000011011000011100001001001100000000000000000010101010000001001000011000000001010011000001000000000000000100010010001000000000001101000000010111011100000111100000000000011110010000000100100000011000000001100000000101100010001011101000010000010100100000110000101000000010110000000000000001000111000100110100100000000100000000011100000000001011010000011010000000000100100000000001000000000111111010001010100101100000101000000001100000000100101100000111000111000000010000000001000000101000100000010100000010101101001110001111100011100000000000100001000000001000000000001110000001001110001100000100000000000000010000000100001010000100000100000000000000000101011000000000000001010000010000100101000000110000000000001100101000000010111000111011000001101000000010111100100010000010000000000000100100011000000111110001111000000000000001000000001100010010000000000000011100000000000001000001100000000000000001000000000001000001010010000100010100000000000000000000011001100001100000000000000000000010000001000101000000000000010000000000110010000000110000000010000000001111000000000110000010000000111100000000000100000110000011000000000010100000010000110000000001000101010000010000000100110000000000000000001001000000000001000001011111011100000000000000010001000000000000010111000000100101000000000000000001100000000100000000000000000100110000001000111100111101100111000001011001100000000111101001110101001101000100010000000000000001000000011000100000100100000010000000100000011110000000100000000000100010000010100100100000000000000000000110100000001000000100010000000011000000000110000011001000101010100000010101001010000011000000000011100001001011110000101111001010101101000101000010111100000100010110000000000001101000000000001000001101000000100000000001000111100110100000000000001000000001010000100011100010100000001101000001011010000000000000011010010001011000110100101100000110000001000001000001000100100010000000011010100100100000011110001000000000001100011000011110000110000100010001001010100000000000000000011000100100100000010101110000000001100101001110010111000000000000000100000000101100000011111000010000011000010010100000001000000111000001001101100101101000010000000000111110000000000000011000001000000000000000010101000001000000011100001000000000011000000110000100010110100000000100011010000001010010110010000000101100000101000001000000100000000010000001011100000101001000000001110011110100000110000111100000011100001000001101010100000110000111111000000010100000010001010101010100000100000000001000100000001100100000011000000000000000000000010000001101100011001100001000000000000100000010011111100001010110001100010110001011101010111000000000000001100001100110000000000000001100000100000001000101100011000000101111010110000000000011000100000010000000001010000100000010000011000100000011000000000001001111010000000000001011101100100000001100000000010100001000000000100000000010000001100000000010000000010101000000001011000000111001001110110000000010011100100000001000110110000001000000000100010000000000000101100000000001010000101010010100000000000000000100000000111010001110011001101001000000000010001110000100001001000001001101101000000111100000000000000101000100010000110000000100101001000000001000101010000001000000000000111000111000100100100010000001010010000000011010111000010000101011100100000000100010000000000100100000001101110000000100001100000000000000010000010000101000001011000101100000001101100001011000100000001001010111101001000000100000110000011000101100100010000000000000100000010000000000000000000000001001000101001111100001000000011000000000010011000000010000000000000010000000000010000001000001110110000100100010000000010100000000000000000001111100100100000000000001000000010000001000000110010001000000000000010000100000000001000110001010000010000000001100000100100011100010100010100000001001001100000000000000001101101010001100001111010111010100111000010000001101011010000000010000010000000000000011000100000000000000000010000001100000000000110101010000000000000001100000000000000101000000000000001000001110000001100000000000000000000000001010000000000011000000000000010001010001110010000000000000000010100000000001000111110000000001000000000010000010100110110100000000100010011110000000110000010001000100010010100000000100000001010010001011000000000001100000000111000100010100000101010000000100110100010100100000000001001011100001111000101001010000000000001000000100010001110000000000010010110000000111001111101001101101001011000000000000110100000000110000000011011000000000001000100001100100100000011100001100000011011000000000001000110000010010000010011000100010000000000000110001011100000001101100011110111010011101000010000110100101000000100001010000000001110000101101001001100111100000001100001000000000010000000010010001010000000011110000000000000000001000000011011100000101100000000100100000010000000000000110010000111110000000100100011011101110000000001011100000101001000100000000110100000101000010100100101000000000000000000010000000000000000001111000001101000001000000001000010000100000110000001010011010001010011000000000001100001100100000000110000101011000000000011111000000000000000000010000100100000001000010000100000000000000011110000100000000000001010000111010000110000101100100101110000001101011000000011111000111101100100010000010011000101010001011000000111000001000001010010001010110000000000000111000100100101100110000100011110000000111100100100000000001000010000100110000001000001000000000011000000010000100001000000100101100011000000000000101010000000011010000100001111000110010000000001000010110011000101110100010000010000001000000000100000000111000101110101110000100000101001000000101000001100000000001000010100100100000110000010100000000010001011001000010010011000000001100001001100000000000010010000101001010010000001000000000010111000000100000010100000000001011000100110001100000100011000000001111000011000011000000001100000001000100000000000000110010100010001100000101100000000011010000000000000000000001000001110001110000010100001000000111100010000001000001010010100000000011100101001111010000000001000000000111000001100001001010101100000000000000000000100000001100010000000000000000011000110011000001000101000011000000000001001000011000001000000100110000000000000000000000000011011000000000010000000101000000101100000011010000000010011100000001000000100111111000011100010000000000010100000000100100000001000000000001010000000010000000000110111100000010000000000100101000110010001000000000100010000011010100000011100000000010000000011010000000100100110000000000000011000010001000001000001010000010001011010000000100100000100000110100011000100011110000100100100010101000000100000000010000000000000000000000000000000001100001001000100110011100000000000010010011000100000100000000000100000001000110000100000100000001100100001000000000001110010000001000001000010010111001100000100001110011000000111100000001011000000111101000000000100000110010000000001111011001001100000010000000000010000000000000000000100100000010000100000000000000000110010010000000001000000000011001000011100000100000010100000101010000000000000000100000000011000000000011000000000111001100000000000000010010111111010000000001011000000000000000010000000010000000000000000000000010000101000000010110010000001000000110101011110000001101000100101010000011100000000001100000000100001011000000110000000000010010000000000100010000000101000000000110000110010001001000000000111001000111000010000001110000000000000000100001000000000000000000010000100000000101111011100000000010100001110100000101110000010110000010111100010000000001101100001010110000000001000000000001010110000110011011010000001010010000000000000101001110001000000000000000000000000001010110001100110100001100100000000000110000000000101000001011010110000010000100011100001110000000010000110101111110000000010110000000000000000010000000001000000001010000100000001010001000100000010000010110110001111110100000000000000010000010100000100011000000001000100000000000001000110000110000100100100000001010101111000000000000000100000101100000001011000000100000000001000001001000010100000000000000000000011001110101110000000010100001001000010000000000010000000001000000000000000000000110000010111000000110101111000000100101111110101110110000000111010000001000000001010110000001100000000001010101010000000000001110100000000001000000000001101010100001000000010000000010100110101000001010111010000000001100000000000010000000000010100000000000010001000100110000000010000000000000000000000010100000001000000011100010001000001000100000000001010000111110000000111100000001110101100000000000000001110110000111100100000000000000000001000000000000000000011010000000110101101001100000111000000011000000000000000011100000000001100000001001001000000111101000001100000000100111011000000000000001111110110000000000100000000001100000010100011100001100000000000000100000011111100110100001000010000000011000000011100000000001000101111100100011010100000000100100011000000010010110111110110110000000111000110110100000000000000000100000000000100000010010100011010010001010000010100100010000001000000001000000000000001110000000000000111100000000000001100011100000010000111100110011010000000000000000000101000000000010110000010000100000000001000000000000000000000001000000000011",
	"0000001101001101101110100101000100001001100000100000000001001011111100001001000000000000010001000010110111000000010001101011011000000000100000000010110000010101000000100110110000011111000000010001000000000011111000000100000000111000000100000011000010000000000001011100000001001011001010110000001111100001100111010001110000000000010010001110101000000010000100000000010101000001101001000000001100000000101000000011000001001011001001110010010101000000000100001000110001110000000000000000010000100001000000001110110110110000100000100001100000001111100000001000010000100000100010010000010000000000000000000000000000000000000100111000010000000101000000001010010010010000010100001000100001100000000001100000001000000000100101000000010100111100001010000000000000000100110000000011011000000011011000011100001001101100000000000000000010101010000001001100011010000001010011000001000000000100000100010000001000000000001101000001010111010100000011100000000000011110010000000100100000001000000001100000000101100010001011101000010000010100100000110100101000000010110000000000000001000111110100110100100000000100000001011100000000001011010000011110000000000100100000000001010000000111111010000010100101110000101000000001101000000100100100000111000111010000010000000001000000101000100000010100000000101101001110101111100011100000000000100001000000001000000000001110000001001111001100000110000000000000010000000100001010000100000100000000000000000101011000000000000001010000010000100101000000110000000000001100101000000010111000111011000001101000000000111100100010000010100000000000000100011100000111110001111000000000000001000000001100010010000000000000011100000000000001000001100000010000000001000000000101000001010010000100010100000000000000000000011001110001100000000000000000000010000000000101000000000000010000000000110010000000010000000010000000001111000000000110000010000000111100000000000100000110000011000000000010101000010000110000000000000101010000010000000100110000000000000000001001000000000001000001011111011100000000000000010001000000000000010111000000100101000000000000000001100000000100000000000000000100110000001000111100111101100111000001011001100000000111101001110100001101000100010000000000000001000000011000100000000100000010000000100000011110000000100000000000100010000010100100100000000000000000000110100000001000000000010000000011000000000110000011001000101010100000010101001010000010000000000011100000001011110000101111001010101101000101000011111100000100010111000000000001001000000000001000001101000100100000000001000111100110110000000000001100000001011000100011100010100000001101000001011010000000000000011010010101011000010100101100000110000001000001000001000100000010000000000010100100100000011110001000000000001100011000011110000110000110010001001010100000000000000000011000100000100000010101110000000001100101001111010111000000000000000100010000001100000011111000010000011000010010100000001001000111100001011101100101100100010000000000111110000000000000011000000000000000000000011101000001000000001100001000000000011000000110000100010110101000000100011010100001000010110010000000101100000101000001000000100000000010000001011100000101001100000001110011100100000110000111100000011100001000001101010100000110000111111000000010110000010001010101010100000100000000001000100000001100000000001000000010000000000000010000001101100011001100001000000000000100000010011111100001010110001100010110001011101010111000000000000001100000101110000000000000001100001100000001000101100011000000100111010110000000010011000100000010000000000010000100000011000011000100000000000000000001001111010000000000001011101100100000001100000000010100101000000000100000000010000001100000000000000000010111000000001011000000111000001110110000000010011100100000001000110110000001000000000100010000000000000101100000000001010000101110010100000000100000010100000000111010001110011001101001000000001010001110000100001001000001001001101001000111100000000000000101000100010000110010000110101001000000001000101010000001000000000000111000111010100100100010000000010010001000010010111000010000101011100100000000100010000000000100100000001101110000000100011100000000000000000000010000101000001111000001100000001101100001011000100000001011010111101001000000100000110000011000110100101000000000000000100000000000000000000000000000001011100000001111100001000000111000000000010011100000000000000000000010000000000010000001000001110110000000000010000100010100000000000000000001111100100100000000000001000000010000001000000110010001000000000000010000110000000001000110001010010010000000001100000100100011100010100010100000000001001100000000000000001101101010001100001011010111010100111000010000001101011010000000010000010000000000000011000100001000000000000010000001100000000110110101000000000000000001100000000000000101000000000000001000001110000001100010000000000000000000001010000000000011000000000000010001010001110010000000000000000010100000000001000011110000000000000000000010000010100110110100000110100010011110000000110000000001000000010010100000000100000001010010001011000000000001100000000111000000010100000101010000000100110100010100100000000001001011100001111100001001010000000000000000000000010001110000000000010010110000000111001111101001101101011011000000000000110000000000110000000011011000000000001000100001100100000001011100001100000011011000000000001000010000010010000000011000001010000000000000010001011100010001101100011110111010011101000010100110100101000000100001010001000001110000101101001001100011100000001100001000000000010000000010010011010000000001110000000000000000001000000011011100000101100000000100100000010000000000000110010000111110000000110100011011101110000000001011100000101001000100000000110100000101000010100110101000000000000000000010000000000000000001111000001101000001000000001000010000100000110000001010111010001010001000000000000100000100100100100100000101011000000000011111000000000000000000010000110100000001000010000110000000000000011110000100000000000001010000111010000110000101100100100100000001101011000000011111000111101100100010000011011000101010001011000010110000001000001010010001110110000000000000111000100100101100110000000011110000000111100100100100000001000000000100110000001000001000000000011000000010000100001000000100001100011000000100000101010000000011010000100001101000110010001000001001010110011000100110100010000010000001000000000100000000111000101110101110000100000101001000000101000001100000000001000010100100100000110000010100000000010001011001000010010011000000001100000001100000100000010010000101001010010000001000000000010111000000100000010000000000001010000100110001100001100011000000000111000011000011000000001101000011000100000000000000110010100010001100000001100000000011010000000000000000000001000001110001110000010100001000000111100010000001000001010010100000000011100101001111010000000001000000000111000001100001001010101100000000000000100000000000001101010000000000000000011000110011000001000101000011000000000001001000011000001000000000110000000000000000000000000011011000000000000000000101000000111100000011010100000010011100000001000000100111101000011100010000000000010100000000100100000001000000000001010000000000000000000110111100000010000000000100101000110010001000000000100010000011010100000011100000000010000000001010000000100100110000100000000011000010001000001000000010000010001011010000000000100000100000110101011000100011110000100100000010101000000100000000010000000000000000000000000000000001100001001000100110011100000000000010010010000100000100000001000100000001000110000010000100000001100100001000000000001110010000001000001000010010111001100000100101011011000000111101000001011000000111101000000000110000110010000000001111011001001100000011000000000011000000000000000000100100000010000100000000000000000110010010000000001000000000011001000011100000100000010100000101010000000000000000100000000011000000000111000000000111001100000000000000010010111111110000000001011000000000000000010001000010000000000000000000000010000101000000010110010000001000000010101011110000001101000100111010000011100000000001100000000100001011000000111000000000010000000000000100010000000101000000000110000110010000001000000000111001000111000010000001110000000000000000100001000000000000000000011000100000000101111011100000000010100001110100000101110000000110000010111100010100000000101101001010100000000001000000000001010111000110011011010000000010010000000000000101000110001000000000000000000000000001010110001100110100001110100100000000100000000000101000001011010110000010000100001100001110000000010000110111111110000000010110000000000000000010000000001000000001010000100000000010011000100000010010010110110001111110100000000000000010000010100000100011000000001000100000000000001000110000000000100100100000001010101111000000000000000100000101100000001011000000100000000001000001001001010100000001000000000000011001110101110000000010100001000010010000000000010000000001000100000000000000000110000010111000000110101111000000100101111110101110100000000111010000001000000001010110000001100000000000010101010000000000011110100000000001000000000001101010100001000000010000100010100110101000001010111010000000001100000000000010000010000010100000000000010001000100110000000000000000000000000000000000100000001000000011100010001000011000100000000001000000011110000000111110000001110101100000000000000001110110000111100100000000000001000001100010000000000000011010000100100101101001100000111000000011000000000000000011100000000001000000001001001000000111101000001100000000100111011000000000000011111110110000000000100000000001100000000100011100001100000000000000100000011111100110100001000010000100011000000011100000000001000101111100100011010100000000100100011000000010010110111110110110000000111000110110000000000000000000100000000000100100010010100011010010001010000010100100010000001000000101000000000000001110010000000000111100000000000001100011100000010100011100110011010000000000000000000101001000000010110010010000100000001000000000000000000000000001000000000011",
	"0000001101001101101110100101000100001001100000100000000001001011111100001001000000000000110001000010110111000000010001101011011000000000100000000010110000010101010000100110110000011111000000010000000000000011111010100100000000111000000100000011000010000000000001011100000001001011001010110000001111100001100111010000110000000000010000001110101000000010000000100000010101000000101001000000001100000000101000000011110000001011001001110010010101000000000100001000110001110000000100000000010000100001000000001110110110110000100000100001100000001011100000001000010000000000100010010000010010000000000000000000000000000000000100111000010000000101000000001010010001010001010100000000100001100000000001100000001000000100100001000000000100111100001010000000000000000100110000000011011000000011011000010100001001101100000000000000000010101010000001001100011010000001010011100001100000000100000100010000001000000000001001000000010111011000000011100010000000011110000000000100000100001000000001100000000101100010001001101000010000010100100000110100101000000010110000000000000001000011110000110100100000000100000001011100000000000011010000011110000000000101101000000001010000000011111010000010100101110000101000000000101000000100100100000111000111010000001000000001000000101000100000010100000000100101001110101111100011100000000000100000000000001000000000001110000001001111001100000010000000000000010000000100001010000100000100000000000000000101011000000000000001010000010010100101000000110100000000001100101000000010111000111011000001101000000000111100100010000010100000000000010000011100000111010001111100000000000001000000001100010010000000000000011100000000000000000001100000000000000001000000000101000001010010000100010100000000000000000000011001110001100000000000000000000010000001100101000000000000010000000000110010000000010000000010000000000111000000000110000010000000111100000000000100000110000011000000000010101000010000100000000000000101010000010000000100110000000000000000001001000000000001010001011111011100000000000000010001000000000000000111000000100101000000000000000101100000000100000000000000000000110100001000111100111101100111000001011001100100000111101001110100001101000100010000000000000001000000011000100000000100000010000000100000011110000000110000000000100010000010100100100000000000000000000010100000001000000000010000000011000000000110000011001100101010100000010101001010100010000000000001110000001011110000101111001010101101000101000011111100000100010111000000000001001000000000001000001101000000100000000000000111100110110000000000001000000001011000100011100010100000001101000001011010000001000000011010010101011000010100101100000110000000000001000001000100000010000000000010100000100000011110001000000000001100011100011110000110000110010001011010100000000000000000011000100000100000010100110000000001100101001111010111000000000000000100000000001100000011111000010000011000010010100000001001000111100000011101100101100100010000000000111110000000000000011000000000000000000000010101000001000000001100001000000000011000000010000100110110111000000100011010100001000010110010000000101100000101100001000000000100000010000001011100010100001100000001111011100100000110010111100000011100001100001101010100000110000111111000000010110000000001010101010100000101000000001000100000001100000000001100000010000000000000010000001101100011001100001000000000000100000010011111100001110010001010010110001011101010011000000000000001100000101100000000000000001100001100000001000101100011000000101111010110000000010011000100000010000000000010000100000011000011000000000000000000000001001111010000000000001011101100000000001100000000010100001000000000100000000010000000100000000000000000010111000000001011000000111000001110110000000000011100100000001000110110000001000000000100010000000000000101100000000001010000100110010100000000000000000000000000111010001110011001101000000000001110001110000100001001000001001001101001010011100000000000000101001100010000110010000110101001000000001000101010000001001000000000111000111010100100100010000000010010001000010010111000010000101011100100000000110010000000000000100001001101110000000100011100000000000000000000010000101000001111100001100000001101100001011000100000001011010111101001000000100000110000011000110100101000000000000000000000000000000000000000000000001001100000001111100000000000111000000000010011100000000000000000000010000000000010000000000001110110000000000010000000010100000000000000000001111100100100000000000001000000010000000000000110010001000000000000010000110000000001000110001010010010000000001100000000000011100010100010100100000001001100000000000000001101101010001000001011010111010100111000010000001101011010000000010000010000000000000011100101001000000000000010000001100000000110110101010000000000000001100000000000000101000000000000001000001110000001100010000000000000000000001010000000000011000000000000000001110001110010000000000000000010100000000001000011110000000000000000001010000010100110110110000110100010011110000000110000000001000000010010100000000100000001010010101011100000000001100000000111000100010100010100010000000100110100010100100000000001001011100001111100000001000000000000000000000000000001110000000000010010110000000111001111101001101101011011000000000000110000100000110000000001011000000000001000100001100100000001010100001100000011011000000000001010010000000010000000011000001010000000000000010001011100010001101100011110111010010101000010100110100101000000001001010001000101110000101101101001100011100000001110101000000000000000000000010011010000000001110000000000000010001000000011011100000101100000000000100000000010000000000110000000101100000000110110011011101110000000001011100000101001000100000000110100000001000010100110101000000000000000000011000000000000000001111000001101000001000000001000010000100000110000001010111010001011001000000000000100000100100100000110000101011000000010011111000010000000000000010000110100000001000010000110000000000000011110100000000000000001010000111010010110000101100100100100000001101011000000011111000111101100100010000011011000101010001011000000110000001000001010011001110110000000000000111000100100101100110000000011110000000111100100100100000001010010000100110000001000001000000000011000000010000100001000000100001100011000000100000101010000000011010000100001111000110010000000001001010111011000100110100110000010000001000000000100000000111000101110101110000100000101001000000101000001100000000001100010100100101000110000010100000000010000011001000010010011000000001100000001100000100100010010000101001010010000001000000001010111000000100000010000000000001010000100110001100001100011001000001111000001000011000000001101000001010100000000000000110010100010001100000001100100000011010000000000000000000001000001110001110000010100000000000111100000000001000001010010100000000011100101001111000000000001000000000111010001100001001010001000000000000000100000000000000101010000000000000000011000010001100000000001000011000000000001001000011000001000000000110000000000000000000000000011011000000000000000000001000000111100000011000100000010011100000000000000101111111000011100000000000000010100000010100100000001000000000001010000000001000000000110111100000010000000000100101000110010001000000000100010000011010100000011100000000010000000001010000000100000111000100000000011000010001000001000000010000010000011010000000100100000100000110101011000000011110000100100000010101000000100000000010000000000000000000000000000000001100001001000100110011100000000000010010010000100000100000001000100000001000110000010000100000000100100001000000000001110010000001000001000010010111001100000100101111011000000111101000001011000000101100000000000110000010010000100001111011001001100000011000000000011100001000000010000100100010010000100000000000000000110010010000000001000000000011001000011100010100000010100000101010000000000000000100000000011000000000011000000000101001100000000000000010010111111110000000001011000000000000000010011000010000000000000000000000010000001000010010110010000001000000010101111010000001101000100111010000011100000000001100000000000001011000000111000000000010000000000000100010000000101000000000110000110010000001000000000111001000111000010000001110000000000000000100001000000000000000011011000100000000101111011100000000010100001110100000001110000010010000010111100010100000000101100001010100000000101000000000001010111000110011011010000000010010000000000000101000110000000001000000000000010000001010110001100110100001100100100000000100000000000101000011011010110000000000100011100001110100000010000110111111110000000010110000000010000001010000000011000000001010010100000001011010000100000010010010110110001111110101000000000000010000010101001000011000000001000100000000000000000110000000000100100101000001010101111000000000000000100000101100000000001000000100000000001000001001001010100000000000000000000011001110101110000000010100001000010010000000000010000000001001100000000000000000110000010011000000110100111000000100101111100101110100000000011010000001000000001000110000001100000000000010101010000000000001110100000000001000000000001101010100001000000010000100010100110100000001010111010000000001100000000000000000010000000100000000000010101000100010000000000000000000000000000000010100000001000000011100010001000011000000000000001000000011110000000111110000001110101100000000100000001110110000111100100000000000001000001100010000000000000011010000100010101101001100000111000001011000000000000000011100000000001000000001001001000000111101000001100100000100111011000000000000001111110110000000000101000000001100000000101011100000100000000000000100000011111110010100011000010000100011000000011100000000001000101111100100011010100000000100100011000000010000110111110110110000000111000110110000000000000000000100000000000100100010010100011010010001010000000100100010000001001000101000000000000001110010000000000111100000000000001100001100000010100111110110011010000000000000000000101001000000010010010010000100000000000000000000000000000000001000000000001"
	);  
  	variable actual : testactual := (0,1,2,3,4,5); -- this is an array of what should really be predicted (first test should be predicted as 1, second as 0, etc.)
	variable numtests : integer := 6; --number of test inputs we are using
	variable correct : integer := 0; --counts number of correct predictions
	variable total : integer:= 0; -- counts total number of predictions (i guess this is pointless, we already have number of tests we are running)
  begin
	for i in 0 to numtests-1 loop
    		result <= classification(test(i), testclasses);  -- calls function given a test input and the class HVs
		wait for 10 ns;
		if (result = actual(i)) then --checks if result from that function call is equal to the actual class of the test input
			correct := correct + 1;
			total := total + 1;
		else
			total := total + 1;
		end if;
	end loop;

    	wait for 10 ns;
    wait;
  end process;  
   
end behave;
